��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�+����Rq�����������+�nS�U�F7&���S����"�M ��U���@�˴�5��.� -;P�~�oa|
)k���BЖ�@�o�v�4ߘ<��4�l��D�4Ak���-.b���mC*��D�i�M%��%�k�~&ʳ��0!����nY�qe��3��ck����o��z"��,f�ը��%$���|�;+#�0f�UhOǃ��2刑�Lc�����|��|����Q��Ol�pf��\�4Y�
A�Y�a@��qnNAz�pד��ݮiF�?��'~&{�X�v����H�	���Gʲ���dӤ�>v�� ���K�B�x��X�[#s��W�V��.��f$�n���:Qn��24"M��<48�}[�� �(�5��t�L�6����ئe3Xa�|=�X$nD�H"ď�Vl��⼞=��5��n�Q���6;#٬"I�L���P����/P=�}�㟂���C���?�ZI�r�	5��]%���ē�2FTC�Sh��Ds]鉬�@�0:�?"ܮAۙ�>���?��i+c��$�vf�:��P����LX�Z��+�'��Y�}�G��)��q��ʋ�X�]���ۅЅ�aڴG��i����(ް?	�P9���y�
�����E==6�iS��=م�gU����!��8�د�§���g��d���B�Rx%��E}��8�!-�U��@=�R ��s�/�ǥ�;,'�f��|�<�\W�21u�a���{-��������k�����@b��G�9SK{[O��Y��7�vb���yS�����	�63ǲ�Sr�,B�/�t�(��� bc";W���"-�����?�1\�ؤ'

`�x��4Q.�H����E�l���5��S���kd1��{+Hڔ�խ8�|$�������؄+����)���gn��+砯y���>3T��Xw5ӗ<,�C���   ̰�78ys
7�s�m�MO���_���t�3���d���*�۱�)!܃�9��-�J���.��qkT�*)�
0�Fx����t�g#@p��s���(��ܐ�q��U)ײ�Zƚś�!����qp� }�̚��=EL������`4�"������ޖK�sW���N�"61�@��a��w��Q�߱��u��D�_-x����q��௖�,���&7�a4C��t;L9cM�����Ul�2s�!��p��Ȑ9�Z�P���J�gO�=�+�v� m�aRT�����֕"�"��iĮ��{���K�9a��g��j"��� V�<N�.|(�\F�<X|��0���I�;g�}��>i��
�<������n�Ad;g�`ZP
���j�҂��o���Ѓ����/�@F��=Z���%֒g7\pt�^�ڐ�=��2<���'�����'$-EdS��2b���A��@/{���%�rT=an\���>��3+UюUl��@� F�:�����	�$�'{4���i&���@5]�ߑ�<t�=R�ǟ.�����KƚzT%؊���}
��p9�;��|~etf.��i��=n�4Nmn��.(����F�&Ya�1_9]�2���u���s�?I��t̋��*��{�h�Ҫ�JMAhbF�j�Z~%Yf�k@�(�|';�V�� ĔlP=�x9���?2�|B�V�s�,^\�^��zao�x񦍸�FC����y�X��R����(vf��ǖ���td���eB1CF#�qUO����w���f["�g53h�%Gu+333��J�T����_����Y~����9W{J>@���{K��-G�}s^��O��2X��B�����Sg��p�V"�g��k
Ne$�s-��|�V�K�H���ӊ�{Ao4�{�u�$�S�?���Ψ��� >���ɲ}���0�Z!T�8�NK��[,L����5N�W f����J+���u��m���0$�ele�W۳!n�@LC��S)ع������$�9�+�N��5c������q��Hް?@_�(��8�ĘiBj]֫�m�$���8��hD��;}��k��e�"�7���þ��/�����ac;��N[����~.�vZ��7���k?N,?��$h��
s���5&T�S�,��� :��-O�W�<L3�f����[|�.����%e�s�%cX`��6,U+E�O1��WL�r��+Ҭ����yٌ� a�]��q�:�Jgf�ߛ�ǵ�\ˣ?��.��`��Ss��U+�I4fG��#�b�Z"�x�u-L腘+)�{�M�΢�u�p��X���d6�9@
����";�XZ��>(�C��!����E	�7�1���%����ļ�.pR�PK%9�٭��S��3���vOb�$�)�X�(��.DJ*�2�� ���QB�>�5F\�	��rH�5.I����y������>)hA^��z�&�n�������7t�>�Ό�W0���XI�??����B|Pi��x��u�C�LL���e'h�4��:gO���3��a����sACg�� �Q�P�+�]���9v��@z��pz.�v�Mz���)+A���O8)�d2�Fu�f�]_%X��*r�E�F�#�ϔO�|%�4mN�� �4�i���B��X\�Q�����-�n.�e��A
P�b�x��ךt�Q��3Y��	)��5х�znl���`�+[-΢@�7�]Q`\yg�=�Y����z��NlUg� ��� �İh]q1��~0֟�~�L���JO�P�!�c�����a$3�׃1`YF�CW����!�
}=4��x#CIw>�5}�F/}��5�Gpk��L2?,��Zvu��,��*j:����nme9�`�<K����)���x��Ƌ>_;m�$�NK���C���TEU�.��Ch�wf>�~k���q�pP3 4���m���4�A���r�ٯ�d��G,�����iez[���f�V]��g	�}Y�s����������W�$P���%"������k=�������$a���ie��B0�^���@���К�oEV:��WX@D��l���:�:��Q��5�9+��1[��<�V��߇�qݖ�H�!.i��8Jt�e�VЪ�Pl�q	%���K6����ɲ�Ե���S��$p]��-vpK ��%lZ=��r�ۙ�˧8bż����8Њ?1�Beo��ϲ3�D	�����.��r�������^��Jj�����G���m2n�U�e�_�.i��a�c~��PN%�i멾�Mf�5N�ɯA���XP&���%I�]s[�c�}ES7_Ź}�B�Kĭ �����9��0���D�f4�Y����+�X���B��9���b��_���?��3IxZ�Zʭ	TM�&]�)�#L��*K��O���bg3�G�e�m�@_k]H��@�#[~w@R���h�&Yw(�N`u`HRL��kj���44�qo�G2�=�%N�)���&p�})��`�\!�]�oi /����h*���d%\��d�@�ƆU*	'X���LX��7V=f �&��)
����@�&�8̦D�&�0��������u�eδ�X�:	*�$���#+���m�5Q���Q;jb��ꑦL�ڎ
`�T�pc�cc�1�G��e���i�,�潟M��[�X���J?t�۹
�>hRT���l˒�}��R��Vj�7���2m� ���a��Y>���T�n}1�H�����B�9�3O�;?z��yi��p�ƓG a�֚�5 >�[�+x���`Q+<;Cۭr�o����+i!��6͟���"^�Em��G-��9�ᴚi�dn�Po��+Y5<>�ѩ���X�HSe���t���+�Ɵ�ޫ��\�~�g�=s�[�%[���<�. ��in-X�t�!��m���"��V<����'T^Е��igǋ���W��pJ( ���QW%z����(��_��H�^�Ht7>�D��)��Ғ��f�n/���hy$�p��c���"n���Oo1{Mo���Tε�j��H	�H��p�΅��5s^G�{�*�=����Vd����U�eX�q��T�x���'x�������g����4s����ؼ�c��w�Y^���j���8 {�|�޲ѫ� }���& }$#�E�U*�
�u
��tA����ޥ�㚶rZ#�hݮ�X�;n����YR�e��H@ V��]�$W�/\�O���) @
g�����r+;pCM�E����:��C���y;���G��i��NW�`ܜn���]�v �����')�h�ܩ����nv��y���ah��ݏ��L|}���`���i��^�:��N\DCs X[�m���#� �O�����������r��@��g�� �e��`	7�ރӅ)��z�:;эjaח��㮈xgv�4�.��b�5.��p����D�~�ݶw<�_&���pS���l���%�2v�	������70�1C��� TJ�����Q#�Dn���B��Jq�!XGA�yR)u�@Z�Q8��M��;��i_k�$��쟷���i�1�I�2�B�b�د��V)��+Ր�z}��q.��t����7�����⢇�¯�ppE�Z9i���Ш�Ƃ���@�c�t�$�CGU�VLK����!ﭶ���T���zW}�$����VM�Z7��N�^�*Ō��
(�'�1���@�"�����#A��o��2'%�j���*��v"���T*Y�f��0^��E&ݱHKT
Ă��=Ry2�����$h��~4f�����D��\�>K!nM$�����sw����W4��;��̰�Oި9Ӳ��j����l�IY
�xFo��˄(�]��������c��#�n��?*İg��#���#�� -�T�����������W�$������z�i\��Ts�5���3���M�JW�Kw뭂�G��{��1Bh�VK��W,�1H?]$ܯYf�
։��Ak��\��pd&Z��%�M��2�k�o/��l�W�/Um3�FdOx4��[�h2�&K԰	.}�q�{E@��!8�������y�������F�0�	�RW,]C��l���c�;��3�/�Yn�+�e�p]�z��Ƹ��� &s�\��8��F�����\o*�'ѷ�(+Ȋ��8����g��`[l�7�+n4M�/�F�/-d*UϦ���G?DS�L��\�	|,/s�e�Y'b-)*���Ǵ���V�G-�n�3et���dce[d�d�Ȟ�j�	���y�6�?@�j >��X�0R���;��C�C���d�8��C�S����$d�2��g��jyL��C���V�k�R9�:���A_�B)]f^�w�O;CСc�A��z�� S�c"�.�0����;\X3�͖r�ٷ{�ui$U_�iQk=�T��I���J%��O��T�rp���i;=�M��f����c����I�������
�*CX�iˌ>"��V�f@bW�������lz
0�+�n�$
iC^D��p���9�Hd��e��n,��J����z�*5A�k��^䔦.�Q���D��]���@�_�2��N?u<\��	��̆��b;W�%�=\��TD1 %K�)3,h�a�.2~��']��}Sul�0�3�̾���ߋVUwo+O*����p)e�<X�;L�>b�����_fg?%յ�B�H����ҧ�	l~�8�D6�'�1]��BlU�*C.D���y��vxN�Í_�<f�[�5ɉz��_���G��c���n��;��yk>,1��C���ɉ��/z���%+��?�?��a���[#Y#�7�a$��l١v��R�#���Y�l��#nN�^���<��X��\p?j�1�ԏu{2X��L���H��;\�
!�AX���� ];�����ւ,4x]$pT��k2\�a��!�p=����@�|���fxFZR:��F��%��5�jy�qkj�)}�?3h�0���$�<N�l$3�,����ս����|#�.u�꽘��k��r�u#'����K�:��|@���@R���� �)hVGD�9Q�.	�;s��Ϗ�O\�u�IS:��T�O�P�1�Gl���^��tn�sNJ0��W��م$���X����hk
7���INԌN_v�z#�&���X�%g�.z(�Z�+O-�8�}Q]b�[W�A���jx˿$�\�2��ѷ�������D�Ah)?һl8�x����S��bx#8��Bں.K��9u`}�HV��{^����,�z�1.�,f�j+`�� �bc'���^9�����lMu�(Φ�~�Ti�*���� '���Je�� i�B j���Q���h��j(B��L�j�טr>|�>�
�' �98�*������}{��|�;2��a�QU1�jV��(����qp�nq8���o����e%�Mu2cn��Y�"_�95MW� �L���4QSY �_N�:���ɕי�|����dj�2Q��c��IKǫ��SG래�������n8鞙��HO��r3z¶=I	��u��ҋ�=�=�d���(b�h8��c�?�+�y4$��L��>����ad�U��cD���ÍD��?��� ��"�/�E},�K�4[x|G� ����%u�g�+:6�~���/,T�������(L��}�`p�Uˬ+��v7�2t�C��07�A�pĺ%D�px�*����u6�>�'�"�׉���!�����(Ut~���jb�����0��M5|�r>z�T�9��Z	i��X�Wv�'��J��BB��&G�%Q�?�E�-��Yl	!�$��+
�Rj�k2r�p��|8�9��#2KaEJ[��S/��3T�~K[mT����D)\�7�,�\ɤ����J�{�)X7p�w׆>Рʂ�(1�A�З���}��b�(,"W�R,ԃW�ͳ�f��%Z���(V�fV�Jw�@��M8��G��m�b:7ڼA����^~+���R'P�I){7z�+x�{�������Y����[~�u*�x���M��"R�rv��[^�"����qTI4�I"��3��+}M�콟ɣ=*�u���+%m��}�Y+�$�Nk�vn��2��1��,�uT��#��Օ骜BA[m[#��y��>��I�@������>��:�?O�ڬ���)��
:�+�������=k	Iߣ��o9���}3J��s��a��u�H>�t>��K����3S���%Q��yY�P�)ۀ��9!�M0���(�t���-�tJ�hN���j��i��Z��v�Eq[�p|W�\-?�2�Ǻ�!�!	\V�,�̮��Ӫ�*��$aV���?���]�0�)��3EOU���r��Y�`��+p)Z���%����@��h B��]
�gKC��Iyڀ������ݴ��4V��u����C��q���d�T�G��&��j�z�Ɉm��کN�0찷R���XK���۹�Gvv�h�"���5Eo?{�b����+z|�겸�ZO�3/�Z�M�n)җi�Bo�
<���qG#�Ҋ5�f�E�5�V�e#d�b�1�/EJx�=p5�zE�]N�̺�?� h�ϲǤ{=Ozfn#�3T��;b�&ɐ���׽�KPUQ�p����y �&�O6��o�����G���<"0�� ܩ��K����yo�
u��'v������MТ��!���-@*����D�+�qSL���0U�N�"�GQH���}`�UZ����mV�#�M>���E�P����5O��x�/ks�
ќ��ϙ ׋�0�V�I�؂��?� j	KO����=}E(L��@�vW����XM/�ұ7X��3 �n��já�Fٌl�ZJ����&���3Us5�?D]�i:-��E�@Ov,ȇ�����Z�z�f�3{��r�z*L�e�>H��2m�T&0ye����<h�>hYNmثxx@��;��9�@<������k��f��/���+A������M,�g����.o��q��k/�:��.��ՋC��O?Lj@Yg\�=;����AM	*n�>�п|gv!<7��q �%��;�� X�ɜVRV4��d!�1�Y�M�x(�^��"T=\�o�+�op�ZPw��<�%��X�������F�y4�
�R�s����A�vV�'鰧���Zsd�>��"*(P8�,���9�/=h!�Ѕ)f�c|�^���FP�6��]�hU�Q���VI���IS��F6���ȁ)"({�RG9��k�tO���iE�2哥Pg�%����mmT�W����n��J�����״~�lh�i*o��H���.�O�#cs|�E��$2���/�I;����{h��������"�p���>
�r�����8A�Pn���iX%v����k�Q4�vy΅�R�\6�	�����	yZ�"�<����\��A(Z�6i�J�G�mN$4 Xɾ(�+TǱ���F�y�w⢍��/�%E��� x�РQ����H�4k}.Z�e#�iR�hht�0��Kȴ$@ ֹ����%5J��7�Cl��<4{��)���Y�����x�.������v@��A�u8�Xȧ/�[3$˥�*VTM�hVo�!a"=�~��3Z�z�}����_wwqC,���W�.A���>��Vo�������-�쳺M��>e?=�`A����6�PCx�6,��3g�����<E�0��(�P�y��o�U�`��n�c��\L��\�� $�Q!ȍC.*�$)��6*l��D���n�dT��3a�s�f��_2U�ܥ��쮅0/���+��rw�D��4ݢ�l�5���Il��ɂѓh	z����Q��C7�S��2�Y���4��궏��M��y��!f�2��J����C���hiQ��d��aJhPY��&�
Y�Zȕ������Ülf1Ꞿ�,!�e�ZҞ�n?	eS�~����e/Ƅy|!�@��a�Y��D��e��S8S�U~r5�Wh=<��.�^�!�_H����/m�J�Nf�v�i����u�K�%�A��%�S��1��N���G,aM��d0����f������/�@u�7oQ[pͤ߉GT��aڬ�f<)K�z ���_sPJ�cB��t��X��;M�^�f�=�9����2���:�B�'B��=��>Zǂ���1���!�fGھ���v^<d��o�(A�B(̧b������`�>9C,�Ŀ�I��hh�8���N���"�,���Q����ǊHk��@t���6L�z����9s��j��K����jx����s�Z2S�������Q��Lix<v�i8��v�f���o=̀��9+�Ek^���߷X�֕F����u�[,�9G��Z)�mh,�O����a8�g�?k;�\�M�-��J�Lp�+#N������A,X灁�Aۻ�Z@L�,dG^C#N9h`� ˩����V�#�6b����v�����:%uGvɛxn��S��?T�:�HI	,-i-�s´J�����@��\¬�s��)ށ0<�b?!�ּ��?5��i�`j{8���i\t�k��R��A_T�`�L��k�Ũ�.O��!aA��.Q�d�w��Z�k��6V���9�f���ځЍ��fA�.��4��b�l^g��9���nn�V�Fj {
�����&�OKʿ����R�X�x2�`^����WY !�`���+�h�ml�I��	�Pc^���مt�C�c��$��}���B�Z%B�W�^j7�	��JH��I�J�3��s�<>��Ic�_���w|���p��>�J�Ǵ��|�>5��1M'
c4Z�	�Z��i3����fɩgU�W����m�Aq�T��oP	e���c,XW'�,L�o����u�ܞw��� `}kPz�,X}O��vϿ��Z�I%�>>"�.�cy��0�s~sm�X����ȷo��w�6?���εQ�g,y���b�x�(\)�~Xu`�������2~�O~��F7���7��Lp���%�]�T�Gî̝�;��օBJ��LP�O/�
_��٢�����뻸�|~��N0�G0�,u���܌s
���OO�Uy}��p�G]v7�lRO�S����m*�F��R�W��i�`բ輪ֱi@��G�'oX���c�e$�^)��I��P<��/	�+/�(�g��W�ڐ�d�������(NA�P�$�1��c(bVAr�9�i<ܩ��/
����@�Pʙ�[x
�˜��L]�'�~b�lX��F�$�����؏�Y�R�P ��#c��j+��:�p���r�a��O��(8bz� 'Trl��Oխ�"���΄��9����})C|��``)��']E�b��P?("u5�Ԕ��H����֔L��%�؄�8�X�M�kǲX�0>'J_�0���A�+�Qp
�
)����̔E���55ᚅ�� �)��S-�@��i���i8M��'�}sR%�|����н�6��c�̚�X���:L�)�q}mu�������`�u3�a�YeК�I`���ၿ�M��WQ��e��j/�/�/�tT���!�+K���9��R/��MxlgI5�"����3
ދ����CK��RWS��\s�VS=�*�����ЃY���cӬ�\��X-�����ڣ�Ѱ�Q��R�aya��y�%��)��Ԅ45mdܿ�&<�wF��SӼR6�zp��uL@-����
P:�|=��x�_�O�����U��Kc�զ�P��ۇ`�c�%2hF�,
a�!#���ݔ��[[�ASw�n���;�S.)�m���px��.i
���T��t&+8Z���HWoTt�����T��گ��TM
S�Nk!�əM�ɧ/\��=�
uoM-����)�(�#v�E����3�ؓ�EX������z�m?���E�$`PjևPk['zGW��ސ��@z��g_[[ݱ���5�E�Ȕ�E撟�F�:��!���e���V ����_4J�h����qUw�*����m�gwy��F3ق���)��ی��l_�~O�����h�y
4Z *�Q�Q�V6;9�̊�	��Rܸ���e��}��ی�+�����`7��Y�I�7ja�B��/~8LmY���6|��Ԏw�.���B�:�{���1��m�@K5�]ᣪ�m��+�� �+�(Z�*����7XѸ�/�?�ވ[��`f�W3%������b�f���wcKO8� ��D�B+�Un��'�i��
����%9����q&oR��\p����1��>K��9P���Z�����5������l��b�����7���;/Ԣ������d��C�["�1����{���?��#�pX�I��A��ۧ�S�@O�c˙P��,���F�%5پ
���b.�'�WN�OL/�e�`��Y�1������W��K-��f_��4N$��?�� ��'^���zh�A�L�Ii'���&�F�K�L4k��5�-P��V��P�S��*s���H����nBm*PKۜ~]�J��D�V,6Y��T��ǩm����9� ��}�Y#$�����kxC�!hj��mzZ9��.1�}��/tF�>�W0ݜz�it쑰�y��� �4;�?&�p��(�<�@��`�J�DK"�m��i��|5�@ഺ��B�MC�j,��cͻ������M��1�����Ϧ��5KH����*�t$+��e�)^\N�w=���W�2O��"|��SŚ�|�b�����[7Q�D�VI��bp�"�xY\i���:����b�dT+����8*�OC�mWM�}�l�L�Rs�(��zF� (�(������6� z$�Q3���W7��(�c�����OO���+��G���Bx�?��s<�N�3 bʖ!�i���#�t^�\�LũUW��:b�M�x@�ܼA�[F�>�I<��w�3��b8�� ��Cg�R�TI<�Z�ك�^��?)�t/�.����ƺ(7jCK���+UC͹�|v���}��PL�����L��a"�;'�5��?'�A5�IaC3�#o�LY+OF���~^�"]Q������VB�d !�#hP�y���\94t綋q����hyB���Q�[�DJdh oL�1z�oh��|D.��D����R@%X<�gU���l��iXwlo&`a�I��Q�P\�Re��gzR[��B��'�`0@O��f������H��!�ah0�n=8�OA%8C�[F\�v# y�A%0ܜH�C�m��*q�8���Ǌ�y���g[{!De.���o���XC����B�C"���Ɵj�Y�4��^��l�[�5��Q�hL��� �5Tx#,W��D�R2_�7�g>ΔM�*�vR��h���d;2]�P���t�TJi������%qp�EF�K;�}�3���nd�	��"�H�����pZmL��Bk�X���G��!��%���M��y�տد�ar����vb+�K'V�]#t$���@�;=q�n��shB���� !�P%k�* �I������5�yl���!-=�ȤBr����`��������4k�i�����Xg,[��)=ƦGf�h��:¬ڗ��,x#G���k��;�R��ۆ2�놎�������2 }��W�]��f��=�6�z_@���(�PIВ?�])}�
��"P���\�7H6�Q/��d��z'������5!�><rC���X	�3	gtu�>�:��O*�D,�=h���D&"(�[U�Rm�m���.*�ۘ4r��S�NÚ���4% �������FЇn8�	�3���Ye%�8��e�F�����~�.d���:S�B�}��Q�{�����Vq��`�"�@�/jS�2�Ԗ�c'�����5�1�F(ᖟ�@����n�ϸ��͢4�n�T�Xd�)`I6�H��d�����G�D��ڊ�A�-ޜ�Q.�(���b<N���`�f�_�C�|����J�7<�0OU��}F��FN;W�Y?N8��%/˃����$FS^�j���i-�o�9��yw���B��lj��f<�=��Ѹn�\mZi�V�>�]73���1������s��ZY|���e�K�	�Ux_��gxg׿%�J�(�u���z����Bb��K�W	1޸����x�0�\�z��}�i�0��{�#L���u Ѐz貲�����j�@�!�:�#�9���ݬCNW�@��?������[�G(jp#�Aɳ9�%�B�.,.���~W�40��Be�-�<�,B��K�?�q|��u�@�a�,��1�S���ܑD��؏J͵��%���	��f�6�A�b,�L��T�1���W�U\��=3/MH�	&6a��� ^�ț}C�pof�d!����[
a"��5وK��o=)���=�J��՟�I�(���S�o��r�v�h��C���&Tt"z�r�4DK�'��?�)�Zz}BZ�,E&��j�Ԃ��.�p��ş�(s�߄��2��E& P�hs�H��D�J�X�VF����j<�	"�9�j���.��{�����"���w6�n��q��r�/���e�t��5�\E�y����a�r*�pv��yN�)��_+o��J�U����������3\ǄjX�.,�|�Lv��Fq�a�~�̖��:�9���E�q��#��(QՆ9���s�Q���}gȨ̧����kӣȦ�oH�_gJ�� ����H
�G�����ǼI�3t�#�"C�)��
G}O�s`'�Y.��ur��N�"�ʊljX�P(	�i�&�^����>[d%�S�N&%��r{g�� �)h����]���#���m|]�@S�W#�Q��T�t/#�DR��Ѣ��O����\1��]♷%+yЍ󴁣��l΋�k)X��'�7zJ��u����ƼEKA���gWL^�/}HU�Q��C8������/�L٩�ƺ�D0�W��������t���N������?t�/�u+/�.��\�g�K4����$$) ;A14�W���V7#YRǟ	�� r�m���7����ԧ��1$�ƙ_��'�h����0����ޅ��dTZ:)4̴�FUCBB� +�!h]�7�I��I�2��0�1�E��$��AH���N����q���v^q?��^�-=t���y�C䷻m�:Y"�B�gT�Gu\��jl��n�q��ܳ�3�lE	k��z;�WG���$��N�E*��m�w��]�/�GO�����,4�;�Q%sL7��x�s2e�N����^���3}�vd��?J�󲪹M��[%��A����j>TDi4	�񁋢���D���t.�@9�~���jM=��`f�����bJ�~,n�\�C��
\����<V����5ͬ�QmU�y�5�ݨ��|-'ĕ/(D�������evc��Q)l��7���C��^��).e��~�T�ڟ/̽⬨�����:2H��R(�PA��_�U������X>�
!�ٟ���(%s(�<z�,+��}~&��yaW#}��pT�����P���E'�V��f��RF�1
��c�,�4�Wu	��L����Y���IB��;�s� �)��/����������&�m��+��aِ��?k"w5O��h�l��np��|�u�M'�ע����<Uz����oi�Ȳt3m[3I�mb��T���Fe�F@���P]|��F�`^�8^�aQe� �K&�xC��V����N��C��A�Q.^e�\���G��e�R��7ܰ{�cg�*t ̹&���$����4�[]�K_D���5TrZ�u�K~zf7�q���%�KH,Ӭ�}���B����&��H汙�/i�q�'H��}��+�e|;��+^Tq��Ʊ"1���q\S]"$D冑�UzjGK�%��y9�΍j�3�^�˅�+��v��tC�&k�W�9=��8y=�R�,	�I���v���Q�����J�Y��~�,/)dާ�\`^��f�x�Ml�� �-�e���Třj�}]��v*l>��T�h7S��s[J�������l�z��2̈́}�O3Ha��ǨW�0�!���b�4e(&
� �t���;}���
<�v�>�g��#���i]G���?�D���=�A�٦���x�M��t)A)���ƾ�n����
+�)Yb�\QD�;��7������,KA�ZR����>.1��}C��*�x8��k�Wo�`N+�m��f٘Rn�R�g3�����jI�����ߗ��[������gxa-R>�X%�o�f�!�n��8��U�&��]��QEm3/VeS3x�7G�d�wIQ�݄*>c��L�6��U__$(~����i�B�W2�S�/t	����Q��c=�j�IUΟ�+",j �px�>�������c��z�wi;�R̋��F��"�aئM��T�d�^z	�����qM����o�{+"�������0#8βj�$�$N�0���I���x�(�
��x���pgV��Ӛ�D��1X��N���/Q����!�j�u�˧*`>�����9�)`s�G��I�T�����9�{j"���O��UWV�0*��E�L�� ��,��U�x���e�-s��դ9�.�����e���Y����7QI!��҄(�J��Wו0U�NaG�<٨���;|���A��ýtAP�(�M�T2��@Ȏ��@��(���Z�|^T�ұ�B�\>g��1em���\?�%���E��oE��ڱ��QO��^C��+�_?3g��ǽ���M'*�J��y̺y���|�*��%*�9�ׇՅ1r�g]C�� ���U��@�����[���0/���U���� ����p��uƬX���gࠁ���Gai	��������U5뤦D �0��p��]^^�f�C~�(��L�����F`��g��XZrf{s}M��Z��iD<����Ԋ�{��r�
��s����~b�/E�,"�}:���eՌ���&�ڑ��\I��=ܫ��h|j��7& ���[�z��������/W#E7��&�0�m�1
˨�w�t0���.��U5�#o��Z�yz!M4�mdǶ$|2���,���&ق|�P�,2��d��V��5tӐ\����{~���t5��~��W_���[6��| Ru�-9n8�v�s'Af|$7�W��KtC��uɯB-�#T���v�4[����dо�ŐK����b�6�ͦ�(����U�5��^�C��8�ZO�8����t�ƕò��Ո6
~`�y�bh�R����R���O��#F�C����g��lw?f���Z�?��k2�y�!��swJ�!/ӭB �ɧ^9�Y�>e��:k�/�w�m��*��酁�0
��&�����}4�GcP�2���wj�IJ -���+�� ��\aYM�9���d�]�*ۭJ������jc��{gɷ�b�^s	TѰ�]�N�Ԏ�!(=�v�)N�uvĎ%eL���1�5�4/�B��0k�k�4E%�&.�z����`��� S֡�+öh���I��	�y����ڔ0M�K  ��9?^b�M2�P�a�Lc��v�t�Aae�ۧ��诮j���8�Ax�х�1ZX��).7�v��'$_��:\�����7�n�C�ǥ�������R�N��2��F�m�C�k.F7>�cȔ)p�$��+����kW2׶L?����T������&m�e�>\C��Lg}�q���<w�~�S�!}�r[��F�%'PUl �޾�c�@���R�'��6����L����7U'��[\#Ƹ(�q�g�a����	������3IѡJƫ�]�a��e{� ��3��` +����1߷W˛��"QŜzz��FsL�G%��6A�b�m�w�����L$����E�j-��ȨT�q�M
���ܝt��gf�G���9ο';8��L�Y����(2���q�D���Q2	�
V/�lad�Eߜ�JaIz���N��l0{�����rhg&�P����F�0���Wp�Ƥ�,JҴ�U&�5Ȧ��ym�7�\]�c�
J��
D!5^�a$�㸵���D��3�X��|��T�D�|�Nu*vOS=S���s�8|��Ԧ�_� +:RAOI�
h���L����r���q}���_�" 39�5T4+_���r�0����G~�H�$���d�C��L)��f^6�g�89����~ۀf��h04�9�*��l5]}H���ʥ����"^��}�e1�����mNA���b3h�	�@H O���O�nw��I�	|{eBX������
���G�Ƶt�fl��NmWt�>�	k�ȜDə�3�ec�4��GV�ðd�S��Dk0�;��텂�-+m�u|�Ȉ���Q�� �R���+�5���eT�b�	)�O)� � ����!3�%d�zI��{�9vC��Kd[�v:ft��ȶ+2��?te"�Șq�9H�i㪔���B���{M�ߨ6M�|l�K����P����i&�p�\��`��gַX��䒇�#�%I ���r_�f�o 5=�A�k<����9?e��L��\�}�7<��pdM�~�4Z^UqO���i�.?���g7T'J�_�#�O<T�6R�Nf�׋?z=4MC�7$�]J	��i�r4��Fa��s�ٵ:ڦ`�|��0���0s��<Na���5]Jl�_*���O�uD/��KQ;Ȳ������V�B�^�;0N�����q�B�p�=����)�	�(�!�sGWD�u�ķW�g�p���5�g."�(�%}�E��m�?
�
�/tO��i.7�CeI���\9���~����K�@�M�C��e8='55�-�o�|�g��?��#,*�o�����Z3e�J	��.7�~�hRY=ʼ�4R'��G&;�A�c��Er�Z�f�&�0�����S6|q��۳��T-��'����dbˇ,��.�������%�i�㵫�͚#�Z.mղ��˽�YAc����*�f��w�I�V�L�T/ʜ�۶�6�x,�ѧvYH5C]��p��dY��N����"�O<���gB�g�0���cs�8����v�x�&�M�/�e�Dޫd/����c�rO%I���B3�)nء�#'"�y�0%�®H
�t��V4Q�z����*&'�o����ǐ㿤S����&;î���Bi���U�+�e�{�J����7��j�W����>����O�����Df�U���Ͼ�s���=)@^��T�Z�E���	�y��[���Nu]uü���W�B[���Ы�"L^�k��v�d����ƹ�&�f�㇈��A�]���ȱ��3��%˛��"��8�>'n��?x���P1���=���Sm��<<���r��n�9�n��|�Y��R�KHS����S�ִ�����0f�M�SÌ��F�TSؒ���`��B�'��O<,���dj\�Y�P��>P!&��p>�}{�~��P��]� b��PQ0�R����" �Nџ�a��T>�[tN�ܦ✂�7�5���/����J+�Zߞ�P���j�����J�Yi����Ћ�D�<�ר?	�ꕥ_�Pw�ȗ[��o�w�e�[�;�dp8�WJ �e���Q���ؒF��AG\k!O�9*��DK�VT`�k�F���Pb5�n�K���)�W:T�Ώ�uM��e3���m�S�"�ױ�|��1���^#� �&v<Ͽ:?�`���B�x�E�x6��J��K�>=��U��Lm�j_�7�s��:��\�%���t��k?/��^��-����C_�N�Q� "]�I �fc�@�|�@��:�r���SF�L*#K�acX]�Uyy�v\�>�Q��E��)�m#��+	�(.W������8G�����w�Q:�^1qK���j������?!�
�����P��Z!�K2��+惃)�wC����x������W�>|�8�7���%m�:�m�Rd4�c�sx"�,x<� �#�ɠ�B؍.��͒��W#�Z���ֿ>)��.��v&�E�hnQl��V�lH�̽���,�+���|"��!3�}$�������}�;`"�eV�Xk����H$z���eO�Z���	��|}=x�
�. �1�nU���#F��I@�(���3��~�2�q���\�>�t��l'��x-�1�Ӆ	`���5�⾺Y��ȭ�-
�'�)�B6G ds���a/��ɍ%+�K��h����NO4f6���v�$��]-[�>t]*^�G���VQj�Ҿ�d$�����l�A��M��Q���Ta ;v�ث6e�
|����ca�-�zфe��WU�ɘ��qu�K���*14��2��u���Mx��2�:�I^4(��t�m�f�/��*�{tP:�,�R�RI]���A!�U���BLC�=�矆�߀��lC+�����ן<����
��mKpO�o��^���Nɖ[J6i������L���˺yX�eL�N�ʤ�4b�ː�e�� ىe��g���at��_����������am�L�S������ݭ�:r�TP��[��魳�G��͋7��XZ�c�n��A���Q򄛭׋�:��G��Ѫ�<�ڢ�4=P��\��]�5� �TQ��SwK�FT_-)+G�ɧ���w���%倠�n�,�2�9�hz��!1g���ƐT���9��qBq+$��>��2VƢy,��HOv�k��~c����N4��{�s��ҊDuk�5[ �H��S
c���7I��� L��*=%��y] ν�.С�i��H`�(d�0l���g����T=�.���|��4%�9t����\�y��_�_�Д����DBaW��i>!�Q�D_5m�;Y��o���}���ϥ2Ĥ�7�@�����͛�
Ck�n��#�JdEb�E�p��.�uh��	�5R����;6M�s�Ɉ4A�VCv������|��v��HC����Bx��o����������0V,ڰ�I6r��:�+�_U'����#T�؁�P��>u�u�к.�R1��j#���s��'2d���o�(%��V��Џ��#y�Q�q\g<&��1-?�˘�����
bq�8p�ɓ�d�ԩQ�'�=^~/bg����fo�^��=T�˙GMA��.�V`�f��L[�==e@�aH�œ�F�D���-���v��8���?�	�pc���� оG�"�NT�t�L��4�S4
�k�Nˬ}P�����J��}/�׭� ��:��칧�BQ�7�`����*Yu1숌�=t�So�J���x��8<���jJnKoa�c*U�y �/���/O�%���R�XhnF�~k����N f%��J;x��*?����\�f&����g�Cۂt�"��;����Us����ȍ�Ԫ��I���W�-�������CW!�Cۜ�CQ���),5إC�~�a�J�5[CU׀����c?�e-��}A�Fθ��Л�]Jݯ�Y���W�2�@�2V��Q��Uy:`lh���`ʵ$��V���F��h�dr8�W��e[M�L��r?U��hS$#(OL�Z]�i�qHp���� �yr\��k${6���Ss�Ax�1穛A�[��
�Z�f,��E����W�j�g'��(8�+����ߖL�w�ݻ�h"�M��<Љ.��s����E,�A��J0�cTKI�����ᑸ�`	��QUy�o"�9�>��Щ��Xd�~����"'��YԣK�_�S�(��)e��{�"l9�w�y�Q�Ja!��vU������y;��Dz)��9q��&���%}v���c�K;|A�-J���o!��Z���gqq��%p�E_�����!���E���%�U	fa�����pł��+� u/cZ�Y�qh�~S:�PzP�t��R���z���%��[:������-
3Ҭ��V���vG\��{�购�D\���������%~m��ϡN'Ř��C��$��+��06XG���=M�yi�%�^<ߓ9�����W�s
E'Hpd!ۀq�V����������O<�:������|wո��\H�Е�n����m��������^bʡ`Q�h�E#L}�Z�¨��XgWu6t��Nu�r��o: 't�{y��Ә�^�b�^U�O.-����+��#nBo�1�W�P���l��nG%��5��"����ը��.H9��&8o�jÁ�Ԋ��v,��ř��7��a8�N3��ڎ/r^Ó)�_�D^Q��j:�������m$��4��O:��E�b����0�O�^,[��g�U�p���#�~����hhp���=�r��LJJ�<BF�o�,�V�l�}����N7�7应�@Q,���<�]��t���ԑ�{�+KDjÚ���a�2ɩ�4�ɶ��]���}�
�)�XmJ�o���%�a�L*?��:�C i�!�ۭ1X���/��w�b�A�|a�|.A��9tP#�W38������ڟ�i?�G���n��U��@��,0G�����K=��&�r+�l����Y���/�R�i��g}�-���5��I��oq��^L��z�W(���W_����f}ʮÜo<%V�t�鏠h�ۯ�/ׄ��{k�(�<!�@)�H]Rʹ��L���zJ�Br����u$(��k�d��Ldem�I�䢰���|Ցy�.cŨm��ڰ�G�,��%�����X6z�2ÓD�/��..�8�,�T�2b0�@��@�8).}e�&l��%��	+]I�4�LClܘ�yV���a��Otݲ����B��	�$������kS�J�Ɇ��/��-0�F�� w�	���7�[��R}�B`�]L�M�#�m�爜5�=7��@��̾5G>/�[`>_=Eۊ���NYt�Pq��a���I52IA���NY_�X��m��U�9�� �O^ρRH��|5�}�C1���Mx�2��Ȣ���O$���]5���Q��o� 8}��ì�F����q	�r��a(�Mf�p���*U�h��㝁[q-r����7:�
��遜u��>{e�q�/5�E��L��" �1ԉ����Ņx~���SW_�(3u��Y�/��ee{���~K=eb�u�"���Ju���V���Y�W�^�#*�|��d�ỗ-K4µ.��YkCv��&�zX7:pr)���x��_���7����֗>��IQ㰓D!��ØW@�{������#�\AH}1���%R�?$T�Ca��x(�xy�����߁���t)��A�PM�:6k2{^��U�d���x��L�� M;��A�X��^f���,	�Yn��� bm(㺊F�Ն����X���r����]���ح�i��T	@Ҧ�K]
�9.t2�!��ðykд���e��C���'�u6!�{r���h��t0��H�-]��ѿαnҏ���X��ͳ�tD�#��>8�,�����_�)f�L��/�����9����_�� !M{�*I0��Փ��hQ78D��?�%79����d]�~������"Ri�՛z�����`�&ty��@/��[4I��m�Q�U8�b�v�cV87YF� �����RA_�
#4`����h��쓛<��0/�Ͼ���4%���XK4U·R����R��4G��EjC��t˓m1��������F���g����AݰŦ  ��dD��H�`�9S�C�D�(�גO�n��k���������^J���2%���m\:nՔ\�B�!;��i�C�8�éջd��5�.\���A<C�_�AWZ��ſl�Y��(}Q}�W°��\x��T��¤��L�u�!�H9�Vi	O�� g��I=;-�t�4X�+q���%.�L7�I����p�i	�5u;:���#<i�j<g��R�)���N��2��_d�2���!����������WU6y�B��?š�\rԢ�Z'�� �Z�J15��粵��x~��f\����Å��G�r���G����3��O�b)�s'<��g�ɀw���C�g&m��%&��e`�'��3T�R���"i�&HMM~��(䙕� �Ȥ��$co�\��+���'� p�|/u�l�6�B��lEG��~/4��jo�i��Q�(��oZ��2�X�	�Bƅ̝��g�*T�J�h�s��I��Dud0C���������*�c"8z���9��� �1ĔGDpE��|j<%��_LX�.7�V�ftT�l�|��l�U���� �� ��[���/���X>q9F��1h	,y�ߡ`�WTI�,��.�~>��2Y�5`�k�]@�����c��B[��L�_%#j��K�ATo�=��=�y�p��b�w-�F-�3jSי�b�G����v�,?W_�ڬ60x�>(t�e����rf?�k'f�"&��i
z���I��Ԅ���9"uq��6�IL*���-D��m�� BI�N[9��ٝ�P�Ҟ�.�O���i��V��ЗIY�1���Mc	����̆k�(=,`�����c���I��R���]R�;�i)BI��e�����AI���M��QD����3�\���i]������s��=��2:����:�W���'�kBMlU�©a�T���,�M-�~=�F��|#��N����T�G�:���K�E;<�배����Qo�����2� �z��1�b��/�@>�1�)�k�jT�/��y����׍5�Z�oG��b_m��+��)��G�P6\RIa7)���ض��ɩ"�Kk���}�P�A�n@}w+��_���^r���<z����1'�KD�3̏��o&�TQM�)��0ו�=Q:���C�>������;���͇�M�_Z��%���pKx�[C���LP��\-7�T
�lҔ��S��c��nH�Mgz�OU�+3���i��Z�#<�^��8%-��0*#C���
�~��¬����e
��YB��x�R���f�k�|�Y
H����(oFJ��N��5��c����P�r�8h2��S��5(�j#�&��
�.��T ='�3He"�H���Q�O�����y�����?4 �����P����$ak�S�j��;%[s_�i����C��f@�M+���vZ.^<���ӰW}�`y̟;ZOd�B�fx�޾��s��1H@�]�ђ�ޓN��Sؙc� ��{�$D!�q��v��Q:Dۑ�d�X��n�O.)W�i�ǖmǄN�%�vbh- P���i�vP�,vE;FI\nIܒ�Γ��|���z�1�ɾZmT�d,���L���z����4�[��=�� {�C0c�����x����Ac�*N\:�- @�sŐ�зOe�N(��d�J��+)�$a3�:��Ke/,尿��֤�-���\O\ǳɨ�Bp�IE�,`]�vd���h���$Ȏe�vϖ,$�Ls*ת��n+v�v�d!�H��Y配�zM�Sgb����0�5�U�:*n\�F"ۡ����q�e���a��+S�t�����j{�	Gvx-,�t�wpv��h�
�/	��N�oBLՏK��l!.�P��X�������t[����
F;`��hk"��~���a����q]�uq�p�u�+k��+Э~Jt��� ��%O�;wȉwȪ�/���s���7^�v�ێ~_P.���,�%~	�e�eV?XV��"��h��^+}���bjM��"E��u9A��a#Jw��g�>�Eͼ�,�:ф��S�:�e�$��/�_J\���`�c�T�xæ�/|�&|�6>�ƀ�^s��X!�R����#�)�)���)�{����;[i���2�o�9�@�NQkeTv�O�˷��]`��j�<K����f$/"��<Ei� Lp��d)vJ��3���q�+������u�`	�"�#�1fV��}n�l�8�A�Ah��
�Y1{z���v�\�O���xk^U*�^�����v�8�	K"�I�>��4�]m��!�s	���!RAq���E������6ﭮ�b��z�A�6����3X�-A,}P�勠q�2���?h�SƇ��	G�`��E�tӂy�95�]Yu5���Z=L|W,5Mij
e�B��.ِ� P������I|�❰��c\��GC�̶��1A:c&��[n���Tk��C�Ò�𕖰�߱��ty#����s����Y
�ô�U��<�ڬ���z�����v�0��|�P�}��j�\x��`��*ܸyړ5JO�罗��*�[���I���ҁ�u)�E�0� ���v���䰯��/�4���Cs�Ă�p�����}�p����O/MK������4��s�+�[�h�H�9$��3hh���
�U
�Ad6��7����,:PkQ8 mB��1S����l(OTo����d��	��OS\Lk�K�4�0�ZeC���$W8l�9.��B����/6���\���(4 ���32��A�(��!_	I'�4Rɢ���1G��sJ�&�sx��m4[NҪ�C�b|��gJ��P�W+�[xh3�{����<���{�S'���P�W'�$������s�mɄ��~|��0M}�M(b}��8v��d�Z~���(?'/��引8�q��~�?���!ܬ�{Vf��	��h�����2���$������%�̹j���R+=z�0Lw��~���{�U5g[;vdԸgsn� ��4���?�v�������de��d&T��[
6��æ��\�=�0��֜����Lͬ8>U�(Nwm� �Z�(� AҴ��k�%��,�І��x��1��:�H��Q#nר�������R�$��s�t�������!�����[�|�9��6:>E�0d�;]}Ϯ�5�ab0lB��P)�V��_Z��R�,�4��� "�zgjXI��<�������Z�I�"Oհ�X.�'��6��~��L�!oF{۵��p�;,��rb.$~�7�|�����Ű����>�.%�z����W4v_\37Y*�:�ct8�x���É���S� a<�p� ��y5��sM	�C�`�K*^6+�mx�ڄ����Cc�_@���ݞ�a�X�\�?4O�'�Q�c�VO�������Z1�U�T�Z�S��M���
�#����T��*A��ݻ�d��B�N��7K�[��ܷ+^�ϬX�k��F*p�K�Cx`}��މ�C�хN8&;Axqu-��Y��2e�WP�V�S �b�3�w1�ƞ(Խ�{ǆ����������	Jk��u-8]
Q\�{�*|�O��t�/�2&�f��&`4���%�AZ�j���M8���AM��kh��i��ͱ�=L�����͗��P1pّx0U��u��� ��iR�-mӾ���ԃ���_�	A�5`dޢ��1.	�w�%��ܤP��Q������EJ���$�~x8��&-ݝ=+�����)ꔗ$k�*��W�v�^��܊s�D����(��H�{�n/*�s�p��W>������
����'�o�п���d$��)��m��y熾OPO( �*=�q1��Z"�if��[�`K	�4ݱ��QlL��woSC���\t�{O8�s��p:�;t"�|���p��K���$���="3,�!Uͧ̀՟�V�"������<*^��|9/Ѫ@�����N�Y�QY$e��*��Gb$K��z��!��g�Q�Z֭ϯXJ(�Ud����������(�����q�@���Ն0�Z5�A�dU��x
�>���ī�}�	��80-���l�
z]���=��������׽��ZZG�"Fqb�kq�Rwԭ�6��TL�r�Z��Ǩ�Ҕr��׃��㨻��?�V@��@Nĩ]C��Qww|�������+tX���X��>�&pW��`Z�T[\Җ��6�(&#���dF��K�
O�1W��D,���]�-xO$͓���V3������l��8�[�_�g"�92%u4��vb�� d;Xj9��;�듇��Iv�"�i�X�26	��V�R(��A�S�b�Lh�L��s�gAD�Y�`
�~��@�EKz��H��z?����U�Fr����ᜒޡ^^oe�|�TD�A
K�.u�?�bGG�	̭�����Dm臝�G"��(���>\��c��.e7�F�P�)	n�}Sۖ��<��Ю�ǽ�_�����,ێFt�������.7t"1Ky���������8��h׽	f�s'�a[��&���=0�Zr�?�|P8��)�3�ǿ��dlC.��̦r.���rB���2a�9}=�4#���ܹ��J��+d��/�{%�)r�ѣ�Oi��kg���\���9�z"m�@5��v�+]˾W]n�G��GsЯ^�=m�/eJ��g����"�z��SZ��G��$+�9���R�׻��(�Ua��?6F��Z�KnX<3/���ꍯ}G��5-n�S x�mxs"Ƨ�R����TΕ'6�n��5k������>kđ�2�&�9�<Y>�*S64l2�M2�Gmt�<Ȥ�kq�O�Ge�~|�ş���_ON�B-��yB_4��9,���w	��fJ��(���Fǭ��B������W�a�%�<�X� )��3��V�-C%~ +���'�,Z����+�m�&�,��9�HK���ӽ��� a*���l�HY�ɝ�2$;a;8��f��H� ���ip	v�ލ¬3�T�����LD���Kv<X�t���i����ͼ�)+}X�
5*����,2u�%p<�	D���M$��Y���`��%�.�^��+����cM�欓&#�Q-���Q�u~~�=*

l���hX�a?و���4��tJh�0 ��"F`/(��A�@��K�2�:������tP�j[�Z&D�Y���߆��e���5!s��1Y���x��	l�f���t�!�E�Ƴ��SO��ʟwJ��:��&d��f��(;����bR�e"p!�Qnp��1(- m�s�o�[��$M� �I}?d��誵��NS[�L2)A������)R�y�9�����o+ 6�QJ���vH�(�䐿��h�_ }Ub���`�P\,=����v�.%97�@㥎�.�\�'���7�d3��c�������Ǻ�<�n��-Jvd��;X��XZ�Ǥp8G�Dy v���<� ��4MD��|���0a�*AΧ�w���1
,?������Z��[��c��l��	Oυ�G{.O����\�bC�y��2��ܾ[�uEx"�4Q��n����+�#^�/Y�@���@o[��}�]�����c�8^r���Im4;+�Z��$Sdv�v�9y.�w*��mo�xb9��y��ja�F�;f����L�?�\�d�F7��\���8�{���>4���@�����3P���1�����)��ז����&S"]����%r����(�q?iI��$�n#���7��G����e���9������oƍF� RQ*K��zg������a��v[SŇ����X���$'"[d�Z[��qڝaC��>!�P�u!�}�b|^�V"&_lm@.���;#�%���g�Bj�Nz��{��1I#~8�?��5�%�(���^��\�Bv�%���J�fWpQ0����>K1��u��̡�O���v̈:.������4������w}�0��.�>����J��&f�XD����Ҕf�����6����;B�^� �ekl�ԚD��\��BӁ��*~��ӛo��&�0.ѿ����3���\��G!oW4� ����֍��1b��<��V[5�qXg�[$�q/H�r]�W� @S�o�/CG�ޏ)5J�<��2�&ѓ��y�'If���^pk����*�~H�^��	�7ج�n՜�h��[��Y0F���=�F���d\���؇�=.\9:�!�A���b�a�,W����*��įMpV�����+��`�*;~C#�8��X�e'�G�]A�Ջu����ۭ�)/���۵�_K�-]�/_�*��fO-�-._���7����k@��}G��.��ۀͮ��_~x�7 ~�t��yv�m��v=�-��Pr}�G�������%��]^�G'L&G���2��x�J�}\���86_����#\9�2m�l��=���I�A�3}�mN}t�-?�o]</��X�$���gB�E�F.;��\;ۓo���Z��W���[U;z�f���<�2N���	����hN��
L#��a�v��Qw�B�Q�d�@e��n�H�k��2|O�&3�L
iϕ�5K+�og�U]�;)q�R
;���2�������/Ǒ�v!�������l=������X۵�j���>�������!�q��l��tҙ/?JEJ�"h5�?�����w������q��*����'s���-|��I���y�C�KD�#;*�TvI�{1\8�d�-�*tiE�ə�+���tj�Fi�`�gp���  F���A{���U��$�Nq�Ӹ�:�%��Xh�D��:��u<c�J|�b����ZQ��m)���F!��y����(�NV�f��&�-���O*��:�����t,�}�Rr-��%YZ�
�5��i[�~�]�{ ����{9M���v�W��d�Xq���PY"��~8se��c��@��_`�K?'J����;n����w��D��o8I1�oO��PY�1xk�F���fu�����7�j��UY�M��^����xE�J`8���I�=7 �eylFk���c%�\% B��hLJ(�t\��y���zf�}�l�m���x�i2���
�δΡ6���b�����s`;M'"�_�w�_ά��֍1����Q�]7�YTPZ�;	^�9b����i��F"F=]@�&�>̪�����&����Pf9�AE3��k/y���KD6��m*�����0?0�Á!�#M8��H;9]y0"	���U��T��6T�b���to0J����yN<��̳
�d��	�����3,/;�s��?�?@��]Ǵϼ���+��6����K?�Y��,f�	�o`�,���v�>[A�x>�# �GT��>Z%�d7�v���4�{±-T�Bv (2�"F��!kd1�}�1��_?`I��d",��3� �CR�3��GϨ��v�w��Ò��^W�L�M��;�(�v%j�1����j|��{������mC��X��	[:8Y�(�8lE|�������*gZۨ�	�8V�p�Qa�S��E�w�G�Ӂ`$
Wk��'�4���\}!�;o�����i�����Y�g*bY�(����}���5�a} �&�03�fP��l;�������+D>:�mQ�>҂��x�{�X�cJ�mK��Q���7]q�<�i򑧰x� ۘ��NĠ���U��:�H[Ω�VL誊�p8X�E�� �̭a�Opf�1�_�u=�w�.�XU�Kk0����/��-�j�6P/��|�F1��ǧ�m_���iF��72<5xꁦ^��S.��	C{)���AY��9��*��ܫ%`_��MR�V�c��Pʤ7�+����K.W
?������j����B88jb?�:�G3�����\���e)�dv1��D��Y����wK"�8��O[$�U�?���)LP��ߩ�\R�}ڶ!4**')��[�98�� �A�wq.�D��3�R��CDp���G/��(�h�:���d6�.��Z�E�W�Rc-����4Ǐ�d�Rg�>�]m�Q�]�����̭�[DR�� /1����J[T��Bw��X;Z2��֥piVw�S0f>�ޣZ!/�X�|Hd �������m�d&"lZ�r\+��k�k���$� ��">����2p��,�8�u�/�F��҅޾6�ݛ�(�7�2+D�n��gf���+��� k|J%~�,Ŝ�4K��׃��}Hg��mfg�F��J��<.���c�����Q��%�g�) ��~����N��5e��т*)/��U4�α��[���WkЈ�8P�ݭ�.�椓k�U�U�A���������{��eڣh�a���#��Ww��jtJLF{H?���ŵ�ی,��?Ti !]��߈�|>���T�f��@�ݺ���r+p]��AZ��� ���+�'M�0VU4��`�����1��.��ƾ0��/8�VU>���X�.��p��S�4m6N�]E��l���?$t>}�W:�
�U�`����C�3b�ŵ��S��}��AKi�'4�i��]��+w�r�9s�s`[:�����E���]�AY-��hjq�'Gn
�=έ(���1AN��]�s�;qT�tu�zLd�L���E]`���aI�(����	8��b��h垲t����H�}��sd��
U(�e�7�ۏ�| @�z3��K
�����ޛٔ�9��pؼ�OY[G/
�,O҅��B;>Vc��gc�t�h�Z=�G��/�Z�JwS�YM\��LtϘ��6x$��#��P��7;˾К���UkZ��+��a�Քp���ݻL�1��pN!ÎXخI�>�Y�
c�t:��'����t�n�5�rK\��'��U��)��Y��/  K ��(Sְ<�&4B�Į�eld��ȗ�L�n��j��`�*�>�.)�^o%�܈��xO��D��p�aÖ��9�g���1\�Hd����I��VN��줦����7��A������`�Y-U^|<��-_�&w������8�5�i�R"��UH�� �{�etݒ�G?��~�&#�S��7dA&�ƴz�\����jL�����B^I!���E���Ưqމn�\_���[��
E��3J1���������[S����������pRˍ)���� Y��������}.k��ް��K��_�ba���s���Ԥ�#�'�����f�9o=5m���ec2�:`>Z2�/��k$,Ҡ�1�%��nKoY(��WW-���s��
#�.��1�&��GЬ\.��8O�f��ߡ�J��!DL&b[Q�="��v�4!xb]�\�~V)[�� ��E���`
�*_[j�o�2��t��1S�N}w���&�kz�T#W%���Sdd����l�����[d`�	�{�⠌�(Pa���R���է~�,"X�S�x��Y�0���K~��Bp	J���C/�G<�=�Ԍy�ǧ*��YZ�����+Cn*�k�B�- 7Y���LD�X3�J�\T�h�_=$�[!�G�S; |�jƝ(30�C�	Tz=�WtN�H��W�<�9���Z��ݍ�P%&�^«j.� /��O_7b���j(��ᵽ}��%6x�����`�&��Qk�d��ij�1�>dy�����tDj4��@q�X{g��'t���`Tk.1�{��`Q�O��l�E�� y���m���C�*�9�uQ��o��\��Iu@��&��7�D� ǀ�(���峻m�qRQ�º� ��yA�)r����}|�`ϫ]6�R���Xa���ꒇ;�;_\�q�pϯ�s�'��d5h����g��15��B$�f<��7��R3�~A
Z*�~����m�9�G�qy)�<i7X��n�C*^�1�H�~F ��!�D�й�pJ�#M���m�!?�Lԧ0�SB��R�D�O������>��B������3O�򳏫+.������~�����\	�=^O���c%��5']l�_+���,�ƒab�,��Ns�.�f��]���y�嗴�L4�����a��s[�k���O�U��7��Cv�H�sP����v���%y/�>�-�Z���;�o_g�����TC���لe�&��U��v�xqeYKVnU[)9m|M0�hXʫ�=���Ϋ��̢B�X���,�����4�s'�����o�J�����a���*���h���FŽ@��T�a��:���}��ұ#آ��%��A�[
�\��"�����}T_��Xg�L[���'ߊ�n0���h�l��0`����X�١أ����l�y�]b�B'�T�6�L�}_�/��ii�_7�7���z/�(�芵��_<o��[!H"e?0��R�<Ɔ��4/�Ȉ���5Y�D���4ڼ=����ρ����n2#2�EqybO�@*���#1����/�SR&���O�^�U����K���� 1��������OzV����T��{&kt"׊iG��w�d�n���ɦ���T4�'f���j}K��������{�%��]
���w�lf���s��x�)e���ʍMghGɼ1������:���v�D\(]PYG���v��������r��p�,�z�E�b����^ ��0ں�V,��@�s��3>�\-n�s�CXMV>��v{S[J�*c�~�m�nF$���{��O Ď�S���9x�J� ��!GA�-mfӆ,;l�/�?H�F�W��C�%ZR������)�0�&���5�Kr�����*Np���՘�'[��G/���)b�^����T*���e �:Uͼ��2</�Y�Q^6q4c�4b��e�>=�z�й��D�U�Hl� �s�����4��؛� ��5�?�lhĀ`�?�J��z�8���%/��y�fq��yfo�%C$���ni�Ob�6��1��D�W�Q%�
�ȷ�+�$񿾐�"�o-hQ��1����,I���cpZU}�X�k��:3���!)�|����-��r�>��3�r�w��7�E%�䏓5��u���'^����XA�0�3|��'\�?�=^�+C�'eӝC��|?�4X�����믐2"olS��[녔_�ocUA�=�;U�h9��ғ���L75�+�m�햑�_�Rt���`n���57���!ڄ$;�
� �� ظ:�W��YIy��F���n��.�(�y����%����F��Bg}V��[������ԕ��:�K�I�7�ZF�;�3=9�H����=˃��}���Q$98H�8���`a���XR&�OA�\,G�k6 =$�x��$᪝�k��*����aZ�{��KN`���';�%f@y���;
���h`�T�3���n��X�l���,i���EK
�8��qB>K�x�A��Al�v�q�%�?Xb�hSI禂��=�CUS����&Ή��J��<�� �z�_���O�MuF��P��5���7��a�����)P��Ɩ���ц��nr����خu����������T����#l�����b���!&�G���X��6�*����9&�y=L�g	����р01)��v?x�����P�4��K3o �'��.�ҫ�~��+��qM��Hk�⁃��	��Q��S/٠(���c��
�և�� j�dW�Mk��"��Q1��P���5�C+��r����3jD�p�~s�=�2� ���x��h����qLE�}n�E��8�0�N����HJ���z#ޓ �$����2h�mN����fNN�W^17z5:�j�5�#�FS<8k�h��3�,�����3v�P0�ǧ+smw����.>�¹Z�����x)�@X]C+�m������醯�6�*��.(����хdLWDRed��4�S�a��>�����������3V�MWi�hS���bؖ�D��[���a �{�VBV\HG���e@����juq<e��Z���<I��-7Ԍ����
}�)پ����t��빲����|�d�5����S��Ƭ�c��3ٸ.����q��a��]����l�:!4��c�"<N�,�f�C�4>rq�W��&>Ǣ�,y����B�C�*���:yw�O�r�rQ�?B�>�ګ�,�	Pc�FQ�3Lf�?�E�M��J��W�ƨ�I_�%�5�~*�Y9��Vȧ)����i(��`��]G�[cc����hq'2��뒚mEǄ�)��z7i�v��Z�fF2��M3]��$�YS�N�l�2,����_�	(�W���g�|�f���q�����f�S��	�br���Φ���V΍a��Q\�떙�i���Weo�p%�_.Ť���ֲ��m�-n�s��d<����g��5˅_�-_��Zᱎ����X(c1�Ҿp�����B7�r���@� �"&�,���ÝE�ƈ��\Fc��~���f�~�փ�f��5Z�,�BZ�H�D@!ՏB�x��f۫ߍrT�e43�]Q+5��o�J�̒X}�Kң��3e�Zwlm�Ī�p�E�DI#��X��-.~�&��ӑ�PEm6n��f�nx�S�
�������eͤc��Kޗ�&�k&P���(���Pr���GB�j�6���ޙ�͞�_�S��`�C�H@��er�F$)4��Юr*�6A�O,<�0]�w�������JtvʱC��M��I�S����o?��3�0�D��&�GCJ�y�����	�`�[�!�U�=���/k��ػ(+���G?L_�L��� +�VF���in!}QF4PA�H<2{��H�?z��J�F}��DK�N��7��˟M'�b���6��Úk�L��fۺ�-y��kcU� g�z֔�9����k���ed\�	?y=P�|���瓦��i#�
�M� N��bsM�T�\���$����I�a/��ĊUۓ�lt)�������|g�á,n����[~�K��z�jp�.���	��o��R"��2��[Å�>��Տ9��+���}����8#&�xd��W�Wu��+��M^VC��-���_)��:��͡��YJ�A��[�r�"� /U�v�ʚ��!����.�����(b�nS�2��k0Kc�S�`��ݝ�uv����30Y'���o�+� �m����n�Ywk�fŰ�F۸
�FC�T�*��1�����#�Ԩ��8u��Lg�4?�s�Z�J�`V��ۺ�S�6�+
�ȝ\�ق��)�ejIa\��-@���/����EJ�VЦ�l����+Uk��	��!�b�T7= AK85Chv�B����"���EoQ(�%P�
3���	��t�n�2;-h=G{�Z�Qp������v���Ne?�w�3WE�6�X�t��<�Q�,��P2�~8�~ы[��>�V�#	r���m�#��!�Y�rj����ק���6P���R	~��q��j����~B�c�Jv��~�G�,,�G�f�?���0l� �ʫ0��fY�n;�3�Zw�E#X@���똏�)5 -o�rK�r��S34~�4��A��ej�]�����؊iQ���ʠ���*����բX��� y�B��5O�cE<:AͶ��s��Z+M{a�l��P���WT_>��ȵ��Ή )oa=���l�i�%q���2����"f`Jկ��K���1B^7�����;�-e5?k#��k��U�36��ӹ���������eX�0���8ht+V@����P�?���j7��(��֦�:�~�;���o�#H������K�=�n+[���:Bz9�6����3ĚQ���#�R���f- ���|�n�m�]<Hpà|ҴՈ�90��S�5e��{r�8�q� i�J�a�u�3�L.��B2�`�f���_�{D�]J���B���1�)��y96$�:��e��T;�Ƭ��Y(,=�:���1��E�7�c���&�[]N�o�������� ��E��.�u_;�L���wIxa�HH���
����4�Z�E&����և-�'=��?���ͻI�a+ֵ�d׈T�c��8�J7"A�7���v���XF�j�uw�^�Z�;܏��4smf�I�,��I�2N�j���#>����y��!���%�F|�r�`�d$��oh����B�d���m�p�1��:�.;#'��|#��l}���V�܏{�W;{��ޒ��\QQ`�[)��3�P�s<���j4�S���E2��<��͐�V����'C'�ײ�M�8��mdR���:׏�T������q�L���v4xEf�0K�Y�Q����2��?}�a"ƾa3��
��j�ft:�<WCQ���t��J��)K{\�4'����B����`����'�f�j���C�%�E�2��ⱄ���Ǳ�ف��XFӪ�Џ�E�����j�#?��l����XI�&X�!.]$`�[()X�E�b J���0c�!l�Y潱�1P��OpyI�1z��Y��e����<;(���)�_�*�\�=-�z#u���9U��#���je�a�T`j#�C@h�G��T&��N��!���8���`*��7�}5 U��l:7H�`JYݺa&�,X�&��7��5P����r
��>2���M�W0�}�	�p���r��"�:�"!k�W���Ԣ?��A�5G���&ZAPv��a�v���+�(/+���c, ����@�(nФ����#i�6H����u�2�W��a�X�M�7a��)+"0
 �w�J�K��5����S䉇��aҾ��Y�6��c�ΈV���ࢼC�a�x�4^���8��&
!I xkf����a�����T�~�]S���<e&�
�uc���ghA/������[�VF.�����Ьj����`@�ln����<�d>ņ囤&�4~i����ar�a�Wڸ��B���xˉ��ڡYd�<�#*dV�4������tؤs��Ɲ*�n޳�O�P8Az�\���h~B��`�#��w #C��������_dؐ��1О�h�:�/N+�GW(�s�#Z��5��p�C�W���#(����3{ef�;�� ��e'}��?X�7m�]6T�ۋ7R��(Jv1K�4��xr(�ܝhq�c:��ʐ���>�͹�x���u���vZi8�a_A���S�ԳhdZ^eq�1h�e-dBC���CA���^5�}�σ�v����6�1v�7�.���5[�^�p��&o�ױ�G�pn�h�`f���H��2�����3���[�V�*r9ԭ*Bn�)����/�y<�������v1t.l���&����
�z"�=`���1Z��'P�mkNz�����#hg�X�2��Q���?D�p�*�i{��"���qd���2�kA���#��)����͋�j�2^�xBcY쪉<�A�mv��WGG�E�����c���G���)&��E*rG\��2<�r�+�#�����Sv�����J�x(�$�g��5|����^r&T>S6L�
�a�^��4����V!�`G����%���:.t~3Oj�ID�W|"�b嬍E�¤y��Jy"!��9�<�d�Y�pE:L<�I{Sq{4m�p�3��:�؇���gevo���N��e�
�Wʭ(S���`���u��,!i7�@#�r���n��O �?�E*�C�,������}���m�S�E\t0C���^Ú7�C�Y�ލ� ����޴��I�y��-P�F	���U�J� �b?��`N|Qɡ!@h�G/���d�,h�D��(������G������q�l�h�eJ�J� �@;쓏Ĩ��K�`�5C�. F�<H��}|�@Ћ�05E ��E�D��c�FoU����nz���)Hאv����;�t�ŵ��ص�P��6������&�!O��u����H$)�}�|�W!I部�*D.9��}�칗&w��q
S�q���۠p��
���
�c��69[�To<����Uʔ*RZ�Ī@�!�ϙ�q���&rx �G
�����daO�x'���n����bL�W��(�|�ಌ�ȣo0|J�[_�0I�g�}���;�H ſ6�op�X�.�ܼɮ��'
��nEI^�g3�f��G]iqi�g�wu�91�c��Q.�r��m8p?�kN�E��&'���F2�jA��=�+����n�|�b�@9%Sî�4H�?���PXl>�3�]w����턖UO �S�l�59A'U&�<�9PJ@5C�%$!�ωml� s�hdB!��I��,W���抋'�m���A�݃}��f�r%̍�SW�3	���H7�{a7�'��h����#*����M�z��l7#6Bu��J~�]���3b���1(H-z����.�Cd��7�FŘ�$>z(��Y��H���:�J����(�Ì������Z=�t��7�%�\��ػJ=�:��i�p��!B�k��r)0���Ę�=w�~����|,�j��8��l/�Y�_@��	֪ ]F_�a���3Mg7L�z�:��ο���I��{@[IWd4��~��\L�k׌@|��Ɯ;er�T�e˹P�����n���H��Fr�/ᤏ��*���u�ȭ��ʏ`@|F��̺1Y��(�E�˽G�����>[GXo����PL�4���e���V1�j�^�\�TC ",Y&��N<�;AdT��ꐧEV����ĸ&�8q��m6#���{/�j�Y��?�Z�$I"Y׿�O2�i�0��)� �����,���6C����r�&`�_~Gߍ޳4��7*��!���T�&S�ﻲR�V��U$�,H%�M���V��':�͗�Kk����,�
_��1��X�aSj�Zy�W����Z\�X�ZGjdXМ��r�W�<�9�q�Ӫ�Q�P����f�y�b�-��+�<
7�0��mSKn�>}�@��=H���x+��H0���X�^EY�CV~Ei�ok���&u(:�Ƃu!T���U��r�uՋ0�!�,���|�>�%�ޏ�-����S�F�3jF��H�䤏�|FI 8���}�B������p0܌N�פ����g���۰~�t�&S�jSp�&�T0+�oMºTM�~���%��_�-�*֫YQ��'�DQ6�
��a�F͞ړ2EJ;F�:9}�w*x�?U�X��~�?�Ca�Dv�tb�%*EiNT�J3GF�������j3Ma�3��!���w �%sź/K�\�<�KG�W��yN��M.�5@j��\E
8�`��,Ě׎g��Q��1tY��t�g7���:
�6��dl�\n��BIПeP���.6�F�Uۚ�4<���B�"in(���(�#��F6��`���<8��kǈ[�@	�	���jp��ys0@����-��)>1��cc�(A�ǩ���OL.�����t��|`2S�d��k���y
m�����>�Aǡ~��ꊦ1e���Yek�v����1L���\�]���L�:�ʎ?��SK2.v��SR�@�������iE�hs�� SL��&����{g� W��z->��g��bI��a�lm��v,��)��M���~i��Gf� �f|!��Zٗ��J�t�U>B����;ĸ�Bh|�zE�7�efM���;�׀v�h1��Wqa���'�g4f�,E�r�ŝ�ǓW@ymq���/�8� ��๼�Z+�.\#!L������3ٷ�z�Q>�<�a�,���e!�65P/`І<Qye��q,���_�+	�܉T~��}[{�����LZPm��M���]���(s��H�h��"M)~rXR!V�O�6�n�������ݓ�6�\#k-蛸x	�(��f���o(���r)�BΫŰ&��q:��'g�۬�0um�[~j/�ѹ��+T-������ڂЩ�$�`�
m$���}γ�ExU���@{�ۍ˟O��
N�6L%�'��h��U���}9|W26Ju���"�8����N����"V �%s����,\э&�q�W�[���܊�ߵ.:z*[y�P��F0Q�`'v�52�z�C?���R��l�
��d=?4��/Zh����O�L�2ח�3#Jחz:��L�tKK89̥]���v�	���hit����H	gJ$o٣�<c(smb��5N����
�ɋ$B���)�^��?d��E%5��P������Eq䨠7�K��Us�d���d?��T&��hu�v,�p��q�"OM�'�><��j3a)%�ƕ���Q�;R�Ոr��k7�e�#MU�?�����F�@_��v���j��39��5�ˍ�����9s�f�@�/�S�/˼�#	�R��Z� ��/�L�͞���*�F�O�(	�:ܛ���r�2���"3D��մ�T=D��#��K�\�:�\*�(�^
�P�iڜx����1�5����!/67 ��ee�H��E�?�V����8�Oh�Kĉ"�}��0_�C&�R�WU���E���s��q�t�Z�	ܭ�b�X�ֲ���^ιrFȟ�.<	8��_�r	ڃ��B�ߩ��v,`b>����^�py�����dex�����Q?����j�^�z;z\�סD��_=h7c�T�^�q/����v*d�v��Os��C�W[7�_��Kt��0¿�_�j��H�\��H��V�>v�~����4ue��=�j�~��բ�E���	�}��"��\��艫r갈�2A�p�,Հ�����^�
��mta�EY��~�R��s��ε�J�%2�/��C�9��H*�U����W��3�G}��cy����o�f��XSG�t��U'Bх��S38�*	�LZ4��~��e,T��ٹ�"�D���:}����;�ӧ����/�G��Λ"u�׺�_�d?Cc	ɀLp��� �v̍�
Q3x���	����S-G�4FX7n���O(H��2ͪ�f�L1��KS���5��;S����E�I��]���@t�[��Vo�>A*����C�|��m��Rx�iJ����1h�nT����v�mV�R�x^Вd�
�Y�ǌ��OF �	���lbD O�P���3�de>��+�u>���}��l�l"���cb��4҄"���ʕaN�G�{X�h|���(o!�T@�IK
j=o���XMp�r�&c��{��O��3����2h��;媻�$es�<Ԕ+�xͅ����B�"Ԅ��h��3�=#��&.0��zA���{3���E�`	��r�P��nV�qʶ����� S�rﵺ�\"z!dg�b��ہ@~=���IeV����@�JV�&fĠ����1�)釢��5U7z�/���M�~�k�S�
��?��4G#E��*s].�_R*r�#Д�������)Ӊ
�jjY��z��X(<�S	�wzt�{sOE܄�,��JM�=dTS�?bG�B�W)���S�>\�Rf�)����K�p�q�@�T՟m+:��K���R�ǔ$(uV�M�p������Ep�;4�c ^C(�6/�+[���TҸ�fG�ʗ�H|{a]0���i/��z�EKҮdm�#�v���ܔ��{�6�����G�Q�<~{�]���@������nV	��Xf&�o{���!�3�hӵ[�*&�����=�3d8v&�(�֜����'2K��R�ʿR�5{�]���x�CW�HF�"jA@����N��� �Vt,�<��e��� b�q��-2n�f���"S�f��S"��ޤ�5'����OJ�g�u��'��~��U*R�?bN��A��ާ�F	�U=�5��ȗ&���h�yL�<v̿\���\�&[��v.��nq��d-p����_���D�����@���s���#s���n�l1��<�7�����A9�����̅^AY �a�\.��5Ӱ&'zColJD��������&��IΆh9�����gR���ch�Y�V f�K�k�d%m,����N4�M��ä����O�;s�?�;��k��C~�~֓PLN܇�7���p���w 	l��M�d�
.{�LK�B�XQ�5\cj��	NP/f6�V8�y��[@�)5j���DP*8�-;��S�ǃ@��7���1��ogD��L�H\���>a
#���1�@���$	gP�~�	�,0�P�u䠀6���]F���f�E�t�4�3˕{���ʤ����l6�6�'�O�뛭�=�9\��G��G�6ӓy�y�a�qK���(�+<�"� �ޯ)T�a��!�3|����33Y�	�0�W,d���;Ԯ5�k�hw���:����. �$r',{��I�Y��v䙸m�J8XY��"k�6�B������WM�U�f��ݎߐww���c�E��D�JH��U�$��7��ի\	|hd�~G��ȏT]�̤�02�&o �#�$b*_֠���9b�z��q=�-$������s��91S�-·}�"k	LG�-����2�(����F�����i �B��-j|�C�\��'��T+,��l���������~��%cG��1	Y�sr�����P^M�Y�U��Ⱥ��yd�y�ɿ]�m�v���D7��濿PJ8E���͜Z��ƕ��x�����^׳�j%ޯ���$���$���i�$ikvA��mƳ)#��s�;�	�[ ��vP�����1�1�tE(��ĵK'g�O��3y�����#��M�y2����Ǻ��0�@���1�q��50�N��B���<��T�j46v1��HO�Tl�Lf�uM�rb���QC�W)d	q��v�x-Ǔ/�Ј0��_-�9NU�kMoO�����hI��&��8�������9�A����|�WK};f���V)?��D!���(��o谅����Q&�c{&ϭ�lP�����^=TY�����%��ui���rz�\-�R����~�sdˣ��r��?#d�፦U�;���7,W�ID����K_o�z��#���.P��(�ɺTXX*�����<U'�q�
?G�R��6A׍C:^����M/F�;��%�J��J�%f�VX��*?f��Q�여�Z���Sy��2�W�?-�ˢѱ$LV�'�go#L��A�\곑)^9�T�+�D�����:��T������;o��َ@n�ӠcvU㜟��g�h�^���d����(�~h�X���߈o��Vk1��g�z)#�M��&0����7���ۦ���E/��6�R�M,e/J̖6t7E(�+�����I�Z�)X��R�~�i���f۬�� y�΁�@��(�4h߄���"2_'C���z����ҹxr���ӵf��e.
_�Xd�����U(�]�A��#�	=)]T߄�_,�:i��3~�!C���q�[W���8Z�k\�����~w�-Ʀ�uB�:�&��R��-#P(��8��9�ɩ:.��?��b��~!Y�J�!�0�4�&�mfb��ڳ����>I����J�Z�S�h�n8�"�ʥ!"�#�H�B�sj���}�/q�	�E��P�g��8�Q��N����R�� �o�wR>�a���_#�1�b�T�:�q�@��+���Y�7�|E_�vlv��6~���Lڹe��x[��0��KC�LFb\�����$x�~�%rZ�IK�ux<��RL� ubZ(x�_I(1�@���:�����\X�DנߕqIS쒫����E�oƘ�ՖK.�)*�AS�_ Y�2	K�͕xc��|��ĹA�+���Y��ÿ6l��G`�-�
jE�8�}���q��$����B���6���ʹ���/(һ���ۚp�w�P���AP�\�l~��;��.oa�$sr4��
��X��K�)a�j@���l89�Kp��ZV?4�m�m����_��D�b*r�.�}g6a����T@���V��ﻚ.���ё��X�@��Oa�5���æfBD�g��{��b���i��{dQ��!�^��"�����K�l*�G������F�
�OO�B�f֐�m��� �wu'6oK��1�o%��!AK���M���6�"�4����GN4(�Z�q�P�݀˕��? �����O�c�ۄ^���{�MYÖ`�R�}�j3?-mH(���~�H;��-�b�yu���	k�y��vJ��G�6`�J��������?��x�ݘ"��f���jg�1�\LZ�(��}��Ǣz)Rth$���|��_!8F�o�*�H�Y��7/�e�B�����/gO��z��l��~�ґ����@@�"���+[��&�%�A}�W (���Tdg�T��ϕ��^�n��$�Ψ����Ry	�
��w�Z0��reb%tU��z�5��'0�	�Q��ܽ�D8����� 풕��DM�=������&�:L@���-G�_�$s����t�j���;�8
�E�2�Ŀ�(�
��G3���	�z���C'zX|�����1�ODq��g� �k�I�y�ˏF��PDq(��-2M�J��hqV+*�_�۵�3���E�y��E�3�:Q��R��+sz��"D�ca��<��W����+?�P#j��şZ�p6�5'3K���:�H36��S"� �x�/�M���I�o�E�A��Y�,�I�6�p]��W�8+�&��&j�� ��U�F ���s��yR��&h����2��[ȑԅ%W�Nm�����g����`f��d��y4�Y�l�}�N����d&��4�3n]l{D�t~1Y6�����,�����R����"b�<s� ������ 7���'�l��m��״ʸ~:%݀֝�a����^�1�T��%���Ե��2����0m���<F���LrX�S�UEp�3d,Zv��a?U���+	u�j���t���×�>�Q���̀Y	�g�?vY<�US{Z
��쿱��{S��=�pw2��`�@[���������#4��')-�g��$m�}/\�~zE��j�o�TA��S��X{<,\��?;!��6�7��&�1BĿ�f}�����(}��:f�!T�嫔�����.?>fk�4�'&f,��x��Uz*��e�n�����풐���#�^�/,YƁ��p�!9Y�E��;	�S.c����B��!�y1A)�^��Juh�wȵސ�H]tׁ�kد��������	�gdN���O�ŕ�m�	x��:C.VC#E?�	{��{��\T�����z#3���/I=tG��jjB�eK������{N��*e'ɾ��S�3t��-�
�?�#��wҨ�j]9��(�>�*pAՀ3˝���k��9i�N:��5���2t��8�^�4r�Z���=��z���v����'�`�Cs��bR @;)3�U�K��qLb��<4T�@`�-�Wu�AH����;n�/��7Q���K(�ڛ0���l�3-���0��'����C�\ߑD�[
���`�ɥ��d��=ۭ4�i��Loٓ�Ѭ_H�J��@��< �g^��`�"wU�7�6��MOj�ab�b=S{՞W�n+:Q�E��I�|_kܕ"�����3v��������
�j�?�..����>��zcB;L�А�á���)C�y�����f�H�_��G��>�u\f��`�F�`��n8NI�<*͞m�Y\���~����c
Ʒ���������t?�S���;�+b}6Ӱ��k���p���TM�@�o��EA��j�z�u���2	����GS	ѵ��?�s���D4Va8����NWV��i�i,���qD���l�FP��]L}��a��Zp��� ����ϖ�>��X�כh1C6\�}�j�<j=`����\D��n̨��+�@� *?��:܆6J�0W�IE�%ͅ.#82C���H�u�
!��&"�5�9�f/�����=�Mw�Iҵ����.�Z̛�(���
���:���h�F+`��0���FS��Y�h}�'Z-�}W�����c�v؞�B��2{��������k���mVu��52,�(���f��O�,�y���3�nq�����A^xI��rg���Eİ�{Jj�X�y�jϼ�V�
%3E�!�a�۞�hu�GHsq��fE
;�nV";W�շ������gn�*�	~p����:߃Qs��<��ď�1�ؼ�;H�G�����4t��՟|��*����w��q����q���h"{���@���I���3�/�U=���2����W��д8<� �
1D��������§I�@ģ�3�����'������,e`G��Ob>�?�6�o&�+�WEB���.��!���� ��]��9V=�?"��<Pdn����攒ks����'�g%ۛ#�X��P�g6!��TR+}�*#53��LU�|��Fp�2"i�u3\�psHŹ���+N��%QA$o��A�3:��*�V�\'�G����&���d���8��%dV'J�2�Y%����n����PFС̳݉
d\�*U����=�UGo�TP�J�B���i�s�1�nΛt��ct����`v��֒�8�?�%0.MF�h�ICڟ�g�tYZ�ہx��֖1���f��V�g�U5龟��c�JI�j�~��c��j���K�gG�ݾI{W\)P���]���\q��J�[����j���rNKH��8c{8-R��n��>[�J*ڡF��zHuw�����(�^-��qe͍�5�vͦ&�D �q��D�mk� f<Vd/��Q��y���x�TC �Eϻ�.�V>���<���J�8wԶEG�A�	!D���$���
8����C����<I9=���؞���t,c��Ò����E)�S��/K3����?�O62�.UP,���\YV_�!n87���B�!D�|j$�-޸�qEDe�e�޲��K�A\���\(]q���&�����姉�َ�������Nq �9b��^�\Hަ�Btf$����:@���-z�J��n�N����G���ٷ�Y��D�`�O��şΏ���m{̙�.E 9����(�X�H���'0Q؍�����^j�p�3D��@#Y>~���(�'Y�W�n�UJˊgW�G�:s�dr�p�7��P��l]'��"l���\+ڕ2b��[}��4D����{S��|�h+�7��gJ��/�ax��Aه�A)��3��C;٩��6 $U�+��	�*t{9��KO��)�wE��/I_����%J��:�j_l��M�Ma����ܱE��d�V��b3�51`�͹�{���2Շ�#B
�W-O66!�!�Z��<��o
�pk��U��Vg���[����nJrƷ1�
	��p)I���51���4�����#�M"���o�W���ܐ�[�n.��J�Օ��+&9qZ>���7`C#�b�����)nf���ղ�L�~Z�{����O�)�,T��c#�oь��R�?b9F?3�a�`�Y���ហ��
��K��q��ÿ�>��SK�C�,�J���Z�)iW��� ��ߑas�~BU'U *|�5�����{��A$O��os�G�L�!�;��>1�7�~#��f˶���,Ҋ(��ɺ�ze:{ʭ�%GU���=�1�`K����#�y~�A�<��!��P��P<��������_��]v���zJŻ��� R;s˪ʞ5��'ѭ@yD ɉ��׼A�5b9v1g������hF����|����q�\�)a�Vl@�˨�_��ZO���]�7Ǹ�`�ܩ�ֵ��%r��}ughM����O������'�e=����>�}ԧG���5�f^w��3-�� �~��A�D<ge�2���bf�Pl��Zv��zm7��LW�u��lh�Q�%�z����0f�
[�!�4:�5@Dz�'��;e�/�Z�G6�^Vx�,�p^��!�S�`K.��񑊐�Q?g*�\tE)�=nb�x�߀���'�tH��
�����pk��Ѡ/
n�}�Xy
��;d���G�:cL���y��/ȒTZwf��O8�x��n����}�Gx]�2��KI���0���)�������U��#�'Y(�۫�u�b0���śڟ寅�: x�pj}T�j�S8����E;xÊl��_���-8|���� L���"���XH�����ox+x��S�A�vY���D��d|]���5�`��&�0�gnwx�l�՞F��⳰���%�B9�z5U��-M��e������'Z�hZ�z�I���(�KfG]Q��N���%��,�<X����Eג~q������6
^���d}a�\T��W1��ˆJ���hS6��޸�VQF�"�3�z��ۿv�#���.V�y�%�;��/<̳� ����q��Y�M�y�{�&�CZ�^,��J��H��jZ��e)���}ќr���[ׁ�°�~	Y<��t6τޢ�%`�]���ηV�ݽ�L-�\h��"֏Vf&of9)i���D���_�tc�]=�J'��ݽY��@��z�d�yqk��rq��0a��Qt&�~��#����%����1�21�ݽQ��2/-Q��������7��!1�#�����ch�Є7og�+�O��m�d���%�f5��_��>Y�Y�.��:�<�y����B'��ءz��_ip_J,�����B/��ϻ�%JuOP~��*$�[�0�P��i�?�D�;��%�H�U�vF9��;,���y<>��	�D��`])���/�{�ä��E���!^��H�����z� N@�_�[]�r6nt��P\5��[�|��u! �~��o�*��)t�`}��0q��I�ڲl�U�?Oz�7f�Kc�lG��0�i
�ydds�W6${��PS���h ���m�UF$��ii����Q���ПO2u!gP�t�����`�3�W�H���� �lFr��/zC�B*�9O�_ϯ(���,G��E%rõ�y�S)(NWG�)	��yiDM����V��<j�]KgrV�$_pp0a卛(A��d�V?��b���b��3їe�}��8��4��AdtY-� m��y$�jgg�s
��T�;�:""Y;=�3L��m���1���J~���mI���	�Ä�ҋ��{�~E��֖�֯�/�pDJP(������P�!n�2EZ��-?Ԃ坈lDl���};U���9����a>Q5�]/(�^��z�� Ч�{�v+��Od���.OF�¢]T(��q�1�zl���բ���ױ/ica�G^(�#n$�`a*�B��
���pI�@�:��-M٭��n$jR,Qf#y�*�:U���U���io�˳�ڹ��M�Y����Zݒm���C1X2uz��� ��R��YX��$<V��j�v�O�ܑߧ�7���JQ��c�2�	�&�q���z���@�T���Bg��-�F��N�h!���E��Ht�Ė�DG�B����XUq6Y��G��!�2��\+�
p�4�M�֝�����O�/}���YR��cVi�POIo�.D������k�����4�u� ׋��謭vV�䶺�r��U�Ɂ��\d�2�Ns���G�4���+�.[���0컰>U�-�L/�՘U��R��h_����V��f��x����<�ǇQ��Q�°b�P�mwa�.U��f���;�P3v�-��c��q�&cܧ&��<�(���p~��	_.��07W�)�UMStR#�,�4(���e���)���!Ϊ���z�|��o�����>�g+�k%�pd���FAF�3۽�u��#�Ur1GF�Mh��>vW�4P�)���E<8*�'��5�gV2��3��Um6�?ip�2F��H:u}��)o�*�P���A����(���{~�#�r��_0�ML��`�ʇ#�m�bp�~�!�9�h�3
w�� �k���Vd)k�uf]���p6?�q��B���J�һ�H+Ssǣ�}r�t7�3���֞ԛ/Sɰ�f���������GNԻp�w�%I/#uL�[z�ѡ�U�z��n�܃^�)���C.���V��� -k���)�=N�*2l+;�_D��]>����vȑ.�V���j֜mM.��ċ.��
\�D�P������4��*i?t����
�f����Z����+�6~�j���^��@�O�EL㉵s5�5A��M��am+�R�b)����d�B�8�y�%�����@�)�U���ѫ?8���/f&�󒉏���RQ%T#n��C��E��R䌻S��[�a��G!yQJǄiC}�
�l-PU����A�@��)c�>� TO�xy	D��{�J����Ps'/XL^������G�]�*�׹���5�Q鉫��.Q��� j.�ّ�G������d���R�~�[�Bk��m|`�G�Q��c������(�obn��������a�Ѣ��F�m�X�h3ی� 3�կ�c6p�Hv��;%��&\!�ɓrzb�������owժ-�-��P�
��jȊ�@��uM)���gb� ��%�1�aO����NR(J�x����^�֩ �G�F����1MY y�+~��r����^ܜe�Qr��1β ��\͟U��L�|��=�����w7�i5�<Y���R;=�	������O�����r��f�r|L��L� �0�i�㨈T��P_���Y��2�A(S���%,Lʗ.�LVT���z��(X d���5;{�X�-7�6�؄:Q"���!>�ĵ�&���"���"k�̠�δCv��p�O�W�(�N]��v��5���mY��oZ�I��^*��5���T����̺>O����t�3N�Yq�0!_�?��ۀHm�T����ۖʊ�&
��;oPN;j�/���$�l�L{]�ݐҟ��rdO;��]x��ւ� ����u+�7�X�&��#��aDJݦ��,�䒝��̥SXG;^rb]ga^5ĕ��
��;��@P�O #�Q��\|�Lt[�g7oF���B�����Qj��%���]z�u�'7� ��.f(���|FO��>���YU��E�^��O���7/��@��9m6N�Y9ȶs�'A{��R@����f����@+A>����l�s|�/ 4ߧ88�U�z��!���o)vt����:����퟇O ^��<��t��/�i��`z�Z���bqV|�Ǻ{��8�"��/RG�&J�	��%&�*���c�5_��WE7�D�!;F>����V�4 �K�ze������|?(�X��a)A���&�;S�J��)׻�zpr�ģ3y�>�z�:-���mɱ�.�-����vC|g$��^{��c��F-S����B�	��M���hK���jv�9	#��n�����uN�*3�iА�i�x�8����DG�F#�R�&2K�����\rw�j�T'd�� 2q�'�۽wk�i73�=BJz����)��,����$�	�#[�5�檶P�2���� �k*���m��De��v�;��?��=���k����1��X}"F�dg��S���IK�3��A���c�欶9���N�s1-y��}W[$��W#p �����>�����Ԗ�e*k��z��
-`�5��썵���>u�W�l�"h־���Ь*IZ�
�����<\8@0]{���������l(�Q3يr����Ě㏯^Am����-��Y�QB��X�q��5��,X��@2.����E��v����1�&I�}f{�����95΃�谓JM������+~��꩎̂W����gKW*wx�gP#�����i��j��5�7XC/�{�t��r�*��(u%`��
b�R�
���ϙ��3�Q��I�����L�`�KC��2��X�EN_��Z�zTt���Qd�.�C��;{�s�7��B��9
p����|zͿ;K�HӤ��;�|z7�l�	����!�:�K=��ze�T� ���#0���eR��4�a<���u�U^��/x��}��&�F_H_v�P
/��@΋1 X�|�դ��[�|WT�K�����6; ��a���c�o�;wN%�P{�2X�F1J1���C���dE+�7�0�.e���x����~Q@�_	w*$�V�4� ��Sw�1&�eZ�����=��$h��Gq�V�ޞ����xK[d�迩Ⰼ[[�q7(���]%�Ʈs��D���xi�ӳ�Ta��F\۽*��=o6�f����r��U��b|{C<%�E�{A��DЬ����Ѐ��(8��q�p�E8���v��:�"�s��<�$#H���=3��\=�"��qF�s!���!q/�*�]Z��a���OD	�è_S;Hi��N���[W���n��op�e��G������H,���xC|--��j��iCz��s�ͧ��5�M^9f֍=�V��b�o��xFD�8E����u����V�09�2&=��^�\.�V׭-��QW�v��&��BKX�ܯ���1��>�N@o_��ןX��'��%m��b夕ݡ�N� �����- Қ�Z�&���Q.�c�yb����	�[�q��!�����D!��#���ē0��,Y<�S�Qpc�7��5��q��F{��?n��V,�(��'�8$C0,�Ky�� <���n�so�d��rN��f(��`:!�d�kx���O)ēXx�m���#vX[��Y����g����)��)��y�*�b,���SH��3��S4 h�UO�/�@I[��/��d
r�"��I�Cs���S),F�����#��n���gAY��'ܾ�<*J�Ng��uGM�1L`��)�ejim��Vv��3�F�ɳ�Z���Y?�	5��"�x��'䥂K�{ŏ�YJ�
��f{������Op��
��yn `�{��@�k?�$�~��,v� ���&-������J�b��JiG�Q�87���T�������TT�	��'@0q񟒧��QY'p�l�Qۤ��qT�>H�Ɂo*@J��U&tK3��s!���T���;PO���އ̈́w��;���ƛ!���<\�$�mP�U���IU���B��9������+�l�����R�����ɱ�^"�sxHq�����0�2�+yДc����3`�a��_�9��@g�,���<D����:$Tk�]�`O�'��2����C;��]��5p�+`�BI�b��̧�GK_]׻�1	��I�����)��n��
�Y�S�a�@�N�&�k�,�����RR�_�~1Pz��L���;a~%@������u�{�`��ƛ�P��X�F�W"S�����E�����F5eڸ㗬s K����7�/Ԏ��n֦�+(�j*�ǥ�0Q�v�'ĕ{�[?���b�����h #�������Y����!Hp���Z��ԇo��)�c)C��M<v�@�{�M ��N�g{���O��޶�D�@�7�)^�8�:�$3cP�̰C�1�s��j�EqE}Sқx�4���:�t���\�q+lL�Y5=�_�V�8�.,�amL(gjm���� ��-[k��h	^����V�q�T����n�W"7
��5���7�;�W�`a�����E�<1䒒5���x����6��EYꂍp�NJ��~Up�̀Ӏ���p��ցS<��v����[?��+��k��6�'�B�4��5��J����Mo�*ߡ�C�]�C`��p&��C�������+��F��d(JQ'�C� ��L�tJ��G Z���~w?�E ��2��YJxi��Q�z��CՋ|5���G�'�����R���/��#(�A�S����F��R��<�6n�ȓ�&�Kw���N$F�� ��_������8kSJ��8��ܞ� w�+�.��n`1��2�5� (��:bd����L����"��#�=�E��N&��sÁ��ny5~��D�BN���Z��܂�#�2�͚w_�{.J�~aTZ�������w���5�`�)���<�M�ٗ�㔮�V8:�� D8�S��	�!+)�Wz[�L��k�S���ű=�o]�4�X���8qى�0�����R��/�pv7q����5���� WA{��!��!���rt�t���Sq��Ӿ��$N�8	�F�޹�Z�p�Z �ʀ�t�4���E�:Vd�
��B�X�R��k��}�wYDa�"ا�G���kSQ�x��qw�}�yg�H;jdb����Pf}��	�rr�g*�*�X�q����. z��,���&@��l�r�Ed^$^,�؀%D.Y�
M���]�3�un�H�!B�P���ë4��e��Z�8=/Ĵ�&�����}�����e�u�^������g;�v��?�P H����:��'x�6>��g:�4�C~'h�+��b `#l���^�]?��J���>4o3�8�L���w��{�#�2+?'����PJn�6]B���ٺ�/���a�oy&�0����$�9CO`C����C�-�'��{+d]�������Ԋ`�A�'�� �ER��C��[��q!�y�IN� ��"�����5���`��ou{vU.&*�t�M��k��Rg�U��f�x���
�_�L��I!��/k$�+�ػ��.�D�h����=�9'�8�m�|�ko:\ �y֤ҁ���M�vX^&6�����I�8��Jֈ�)w5*�����R�r'�tӟ�[\��������q�
�M�Ȓ(���z����d�S�Ff���3�\��T6�zQ˰�⸿���˞������+EeE�z<���	�R۷�Tڟ'���^��r橊����"R��<��Jt^���+/V"CM�:b� C�'���8kt�*�oX�
�3) �=Rھ<GI�o��U�)�x������1"��q����'N?��u�w����I:M$�R�[�y�3CC�#�!��P��Ix�|�w��_�5)V���y]n`y/��(tQ���L�.&wb�SrObo+����d�X02ܠ�s6O����B'�T�)��P�!ş��>�dY�m��(�u�fR�V�.@̍��P9��R%S��k�9�OA�4��&��6�����c��Ub�[,���.�;e+fFM�'��]	�j7}��@�ʔ�F�ݘl�łr� ��D~�5Ƅ{�
��M<9�|g��$F���9h�.�.��,�]�k!�/����Q�����$��4`�q�jE���^��ͥ�3�]�@���NzH}C���#K"��X�k�
��
شoP!Kު�E9U�����]�َ3�\pΰh���0U�#��y��>{�W���8|XD|X�It�k�{�|a_���-�	�i�&�k�܎Xǰ�!�a�h�Dך��I��<~�2\�p�s-GGM�ùq)\G�\�x����o��u��H-X�L��~ۼ=�U������ҞS�ى9rM�0�;�����v���o�:!F���g��O2K?��N�0l��O"�n%#���ۡ(C�#�
������m�$�Ӭ\y=ҥ`�ş.�'r�9&x�Z#���,blO_��R��S
�iȈ(���9���p�,��uNB�Y����C>�N>�^�
����H�� k��ҹ4�!LK�ĶJ7Ψ�g�RU�B�����Uk}�Pv��rڵi<�gĢ��^숩O�퇷�ŉ�e��J��۸�ŗT5���P4�#_m` ���`F��с5v�P�:�	��e�@�h�cIC�f�u�f�yn�}���I��d���K�1�{���zF����ش��ـ�*1N�O���������'�Jߛn;�8�� ���^�)�I�� ����]�c��_n,�f@1>΁�%	�i*�jzty�D�|�aFW	\��j'
��-(\d�^��C�sGu�khU��ϻ�j�·4���#�X\4��`�=��f���Q�?������x&@⸪�Y���8 ӉQ0J�cg�D��$�"bhӮEcf�z)w�(<��Y���i�@#T�j���k��!s6$��Z��Z���E@�tþ��p���**Hzu��-�ټd�b�jV7uw���'��ՊL[��c���s�`��VCXHd�K�����P~�9J��S�gf,����k,fb�J��MO�o�el,�%�����	@��PBr�b�C�|�Ѡ:��� �9[Z=Д����]Й�����Y����6��#1��7�PR��`4לo9�OE��+4�J�6��2�Az�s�%��cL�$\����H���3ϐ�?�\�.���V���h������tC�ٿ��2���N<h��\#Ո����+��li��D������`�!ܕ�M��U3��/	����Dd9,�2iz���O��b��=ñ�]��щ�i���i+�b��دm(��׮Ed���.�1�k
�;r;����Y���������,<��6���_��9��wY�p��䛐6�o�ez9"���=�܄�Ѣ��c�-�N�	���$6&]�,��pE�ֳ��jF�`��x�hB�DE��\��μBl�����JSNm��8Ŵ&�Y�ď�M}��S�X���S^~x@����8ֵ�M:���1Kr��f6��w˕�*�A��}��+Vo\��,�.�����ϰݬ�G�93�]�Z���@�ȫ�n�?���'�rB�@�@���v��k��q�W�ƣ��4+�b�V��p�̴#��|d����ՠr�s��/E�H������3Jz�l�7�Pԍ|��]�>�׮���l�#7K�����%�gjo�����V�g�מB�R�+�ĿA�%�xU@C���?#��A+O)B4A�FP�6��<��'������=�H@I��@��)c�m@ώ`�v���HB��=��
�����y{V@�)֑��k�����ׁ$���@�n��㷶ow��Յ��8y���*� ��=�U��w ��Yz�XP4�����6*��>4�,����d��-R�Vjʌ�˰�F0��A�ƴC���Gm#g�7���ʞ��E�L2&L�j�	�2��=�5j�xv����S.�w�U�KFsF�!K���|E�Z؟�_.:�8����YS�L����7gh$n�?'�O��X�`�s �X_� n1���X&$`p��S�Chq�j�r�E���0�b*4�ړH����g|i������]�SW����d�<��.ُ�����ɡ�����s���ua��ҶHܴ@�ʥ 2[��>�C`B�V��c�p��%��3���
��Lj`}�`n��^��d(lĆ���F���Y�9�r��T�Y��P`D��^��H&Bٞ|�Q�ǃw3����!M,b��� M�M���8��5��3Y�I���+%0�3&�(�{ �Rl�}����-8	ke�K���PN9 ��MgJ}��B�(e�~����P9���ȭ��i�ܞHw��{��0�Q��_x�S�Y�Lb��Bn��r�`)����⸨��yk~�̽�����!��yԑ�H�
3��^�f�d<���b��IG��V����u�6iO�n�zRh�fi�@�L[��夔��ҵz��(�GOL�ޠv �����$�����Ѭ��}��y�b���Z�)f�Az,���'o��KM�m>����_RG;+pC]*��aۯ�*(��
�@��Z�$k&���`��&K�S� \I�y��\��/~1�-�;:���c#/ccm2���Q�a{�Og�?�Qtn�b��Iػ����@�M��o*��a+�Q�%,�R~���%=����ǚ�Szq��S�@�"��,�&�R7�!Z�+�/��c=����G)	dlZ�����ڕ��CW7�����:�ȗȼ9CY���^F&�4�U�C#9�vmVT��xi�͘�(C�����I�6��b����/�}=�p��,�Υm�OփX�~����3�j����W%V�4�1��e�]��^�`�s��\�>}�K&��O��2�[9�.Ђ$�U	�*ȸ���_�m2�f��p���p�M����݄��]&65o��p�/`�~3t����>�|X kR�~�J�5��g@��}�7U?ߏ�݈r)��A0��9�V���D���O��;hK��m���)����;�G"}4w�Q�액ȡ{�;Sj�=����gK���>�=�����\���m	-3"����<S�j���F�CX����]x�Hލ��)V=劾AW8�����olׂ[q@J��� ����mL�N*@��u�U	Q�}�1�pr%����c�G�蓼�K􀥜�bG�4�A���bڼ^rk?�9���
�J��U��@4aS�/T��}'0�iܸ���FP�Ȝi!�q�8��"�놠%f��qb=�1:�҃�{�y(��ptϓu�9xFg�Z����&g9�]�sQ^�˂�� V��Sץ�38c��:'�B@7F��꣨|�ڟz]�(3�,��z�_��t�S��/[�Źꭿ�iў�_\胟w�}�h^���K��%৒��Ȭ��R���O�1���0������v�~Z37�D:�e���LO���E��h�.�R� 3r;:�9���S�"(b�����;�0؊��דL����,�N(|>"���A��`'�uw���P�r0�D���k��q`�4��Y����sJ狗k[�2�-�S�t��Eu��bWs���/;.���_L��\���N��7�Z�9��� �;�ⷱ�_�[����UJ�ڤN/ޖ�,(A���{�Vy���`o9���L��1�i��
�LK���i�d6t�9Yrμj$}���L>V�gl����{+�-J%����M�n�^x�NJ}��a���`x�]�U?�H���^W�-4�����KDy�EF���c[��=��#y�$\��<Wb�vwSR��)�9����z9h:�U�޾�g�;�0~��·#�OUz7u�O�<��:
7�n%bA��4qY>|H�n�0~���p��:Vᗫ܅����A7��!ߗ���НQJ`��U��.�0�f ���{ꅬ� �=�����\O:�쭐w�/��)3�jR��q�t���E�D�U�Հض��ۤ'��G33�^QH����|l��@���S�e�w/���G�,���Ӹġf���W�Z<�������\��(Z�%r��(.���U��
C��ȈJ껵vo�t���ot�<�u�����cȚm���������2'gC�����&-������(}Q��q����B4G���I.ǀ"���/���1~�
*�")J�ڷv�r *��}%���W�ϔN�A|������������&V�{ݥ[����#�o�<t����b�wZ�
"�]�L� {��s�qW����bL�mU}Gax�qq��uՊ���ы���f��oW9Q<-�H�ܡ�~/뀽�'icz�*���D霳�IoNg8x
��@x{B'y��Mh�J�孳4��ȡeY�{�x��-����~\�~���!��K�t�|��Gqpl����r�����gQ�x�\���c�5���=����r�.�`�O�}�8l���z�+z���EP�4}�tRʚ�"�����`�ЬN8��҈�`|S���#L�q�v�~mÑ�]�|���|.F�ν٢����a/R$�8��Sg!��I/�!�@�ܧ0ng�6�V��r<l���;��G����F�i�ˠ M��d�u�פ����N�!�����9��M��L&�ӿ2��iG�5�<�0����x7�!Z܎�B�H�j�ҫ3�`�v���g�5M��O�AA��:�D��K-��q(ͻW1�����N�Tf;��YRU��ۉ%��A�(�zr�������~����I.m���P�;vb{�mV3�0fq�����6��h���b}~Z�6��Kw��ڡ�0)c&��'�!y�I�����s��$
�HN��]�/�t���I����)�W<�T�Mu����C�U$��sO��aj��h�����h����P��ۏ*"l֢>cG��[*
M�h���t~�'^�y��^��.�l����1�U���̀|Ir(�J|�v�S�YQ5!QD4]�)�/��h;�X�b˂{�!"�6�+�0-:w�xm�R8���;�s�x �f+WK:��5�FYCd������� ��<sĺ����^�������ov��Y��+���! �{���2����WW�:'�f��E$컧�f��
�!r��dղ���0�є��!�\]2]v���m�RHlL�?D��Ъ{����	YF��݉�(��1M�`8�{}e��Kg��2���z"�����Qv=�8��
�^�Y��^s�d�[���1��M5`>IK�bQ�8�����c�| ��dȩ�iп7_��H�Q���]U���',�=V��=�.y�V�f6ڹ�m@�U�%.9�n���u�_�j���&[�C�e�Og>��?i��-�#HfĠ����_��Ռ�� �)�
i&h5i��YTi�`�/(�� ߽̻^0li�	zWKǥ:l.&���5���V`F��K~�w�*�i��%��,��	����e��ML�W����P7~b�g~�.���	w������񝤂c�t�LO�!�B4b�O�y��r�~��ͷ�2v
g.�pl��*\ʀsx� �Bl[��'�ׅD�f_�[O����E'p��sW���eӣ�um�H-�ض�i�����l��%~Сs�u��y'���*�˷
;���JLg����J�n�����	NW[��>�#�� �۔A.�sm��A��Ą
)z������+�c�����@%��t�C���Zr�Ԩ\�4��i�d{��|F5�`\C�{�����f!D�a�kK��_Mm��XL=g���W_n}�W���n���Qo�;���r>j��^{c�г4<;0��T`��E̺ǻ�9 �B9�7���#�N����o����Pr�ظ���9��"�"��b���f��-"�����I�{��{��z�l�>y�����{���~m�s�)!}3W��"��Dm{v,]L�w�8Iw�+�h��&�)���	9������O��6r��ڹgO8���M��0���_�����I�������0������apU�ă)�����s�m�tܩ���t���/��]f(�C��k�	�fO�Yh��3I��/�M�I�R᜝�Odryyy�j�$�5���F�m�N%�$ꚲ�W�g���R&��f��?A\��"+������=�&��XӲڧ�L�\.]Ϙ9��m`��މNd&H�$���%���F��j˪�}�.�=����	�Z]-`�}���Jl{ȩ��]���B}�jbԅ������e��*`�|�ϋ�o���.]�o�5���{���Ԝ�;}3�~�	�e�E{�P��3�K���D��@���F����W���5z�n{z��{�0�E��n��pmZ�IT��%��� -����viɣ?������by� cPe��M�}���U��H�[�sI��~r;���7K�0�lK����ps����i�����A "���f�Tĸ:Z~�d>�Q�G�?�\�R	�����M��;%(��0= /7����;e���C2m��B���M���(����&(���ܷk�%�K����}3��"�L�@����4�:��8�,�{$5���q'����OX�lO��B�����]A3��5�Qx����eQ�(��:h�]�ջ�>�(�}��}?f	�~���9mtd΢T�#�`�����f�8 h#[b\>s��ӻ\mI�����&~>�|60��`#����?&����W��Z�)w�Yh����t�J����C��M�Cs�����Lʎ�
5�T��,�I�wymů��݇��]nMa�9ف�I�л76�{#�Oߚ% 7Y�ࢰ(!�z�«�x���o�h�0�~�Rp��E�b7V֓@��vY3���L���F��ޜ]w���h��&��f�U��l^�����ۜt���]Zsbi@����x�`�(}:��y�����+�in��c"���f�?���*̓7�v\����9���R�.���ع/��L�-%c��M6d��d��!fXZ�/��sԍ�V㱲HY,]���Pa���}�z����}Q�YJo��K�|��}�l���TGbr�\t Ynn��	����2���w��_66�����x^o�4��+��J�?YX��'0�[m�It����M�UY
���6��/�3�7P��K'nЎ���N��n%��{ɣ}jN��u��u� E����~�:S�Y�F%���u�V��`�z�T���Y�l�B��F$ѩ̿5��+�<X`W1��,@_���^�h�w��{o��4C��`d�|�\�{!
���a���c�6�w�˫���|86�bc+<A�E���C2p2�s�3质�����z�&i�e��K�;���=��YM�Ya�6ŀ�]8��� q_�l���	H�:�G�i��e�e;夸'D�4X�KBZm2�6%G����|�������ɟ�M��~��"n����uc��Kl$; U������/T�PX�5yٮcQX�X�����!����S��3q��@K+��h5��U�����gJ�'l���bf������-l�`��ʵkvLuy�$>�A[d{?o�/1ER�PP�?$��&uG\Bu'�VI<;�ś�%�8�r���n�]�*[Hx�O($<�(�j�O�k�R�� ��_⸏�^v|s�g����2�7�S�p�=�(���
5����ʠ�@>�̷�Ĩ�&�5�ɠ��Q>������~Έ� �L)$?e� `�����B�O�nүG���`�~`q܅���@iQ_�ؤ���O@�� s�=��@u���GS�28ɬ��i�ݷ�pΪt=�
B���I�j�1mH6����]J�{��|�����L��c%��B��,��]��7rm/�3if>���]u����U�<,�\��� �+��,�L�U����O}�}�Z��\��N��q7C���F�`<i�kj����T(X�y��e�	��l����ƍA��m�ZOi���-��5m�A�ءhL����($q�TH�Qe���fo��?@��P�� �q��̖jƈ���s�����{��	G=��i-���O��QL�w���$C��9��7������NՏ��P\,5h;�ǦnjɩpR�]C �Kt���Z�6�l��ܷ�`�]��Au�֮I�l�����p-�%��1+��$��Zfrl�R���#髮g����W吔�7��<��v��"s������ّ��a� C���
2�����"K�"A�%JX[Y#�Q��"��̿�KXL�l�,e�G�p����'n���S�����Ȱ�ێ���7D�����©  I=����OS]<� �W'׺ŗ�O������94�q�r�\�!�sV}�R ��<x8H�������R���?�[_���hZ�Źcc�����?�no���L�����s�`��5�]b���u�]!ۖ�6\;�b��&�R�i3�,�T��������W�R�wc�[V�w����xLD8�g$����.��T��kҾr����$�k;Kv�y.5}~p�y�0�	㤭�J�Οr�/r5�eg�s�C����z!�#N�{��ɪ�L�*�挺�)O��$��PG�6��%}I�#�0d�~�3ֱ���������-,�w�7E9�FFxEp�����J��,��i��b��v?	OD��Cy��vw�����=Z�@U�;	��f�:Ák�P P�v'Sy JO����;��9l8�]��W�3x���gˬ�x�+��rå$}���7lN���2�=S)���" Q��K���@�P���|L]�u�ZE������~��^N�D�H�V��9���>Pb��uI����H�	���u�s꼩�b���~�}l[I�7/��s�h��)L�ax;r�~Ĥ�7�t�o���q`F�/�U_T���GW��ܚI�) �u����i�nIC�M�����'C��#'u[/mh�dj\���6sB3��_����>�<�$w�0)��^D� {+2���Ɩ� :#)P�������~�s&�����p,^]a0���|l	>��0�"�jz�J�*�:�`�S�'��%8{��I}b�|Ռ<��j$�%��\�K��b�nv��]��X?=>fK��Dt�%�*������Q^���#�Vz�p^�:��n��h���P�o��Ok����;*d��8�oמ}���@q�N��)�*��Q��jT�Bn��x�@�ac6�H�Rn�b�7.��N�Ps^����9�Q�@��������M$I�Lk�1�]e ơ� ����;$�##���ev��Ǫ�W�ㅲM]W��={
�q�KSh$a�K\��j����x	��H*��l}*���s���^�	U��􎟌�uUv�&�'�adkt'T�Y0!�D���Y��#i.N$O ��ꃒ���ǡ2��9�2d��ݨ������τ�x�F�v|�4s;��;�$g��}���q�|����i��I�\j�kv����M5�٩LP�?c��Nͺ��@۶������{.�Ǚ���#�W;�p��p�y/=w��z��00[����+h��Ԇ�c��V'��ђ�Ib��tF:��I��M�>�7�ev�
��/�:���2���ԎF���T���
�����F�A��}ٽȣ����������N߁@��{��;�>�^�
U�~]S���9r�*gP�V��iZ(z%-��{.��̿*; [��|�@;(qs������MPcx96�ޱ���7���'��ZqW'd;��S]�,�-��9�4b:�qFm�#O�7���Cuk"WT9uZ��6��d�G�a�LF����oG�k���o��Y�|�x�4�F(����X���;p1����qE��]���S�F[/#����@���^�P ��� �n�f�����zq���yZ�o;cu��gImyHV�v���虣�$���j[FR/@- ��$[�*�����3J�"������eD�n�#��%�@���:�	��B>�`!�\�N�����F��YC���r}p�.G-�r8�w�)���hl�L�S�i�����g��&�@���谺wF ��bm~X�<^FE��TI}g���lK��rk�:T`~Ж�M>����&����m�4��>g�Z֠��]؞|Ś��u��!~�X|XJ�j��}��#���':��Ԃ#�m��J�e=֯�\`R�CT2�B{���W���z��X��T�݋B���mYe���'�� �4Q�;
#ä�%<ͼ� N�;۝.����W/n= ���t��X�zA$�++=���>�ˮ����L!����(��OC��+��d�Q�a����wv����߻9� _���!�7Xo���������:BE��ɥ�1>��g¬�r�֢�QГ�㎹�����L�C�j�ńvڻLiV�Q�_���+�m9&?S.SQN��>�W��k�v�?I�S�Ȟ�������0{~r�[����q�'{M$+��Y���U�
���]�S���V�:G�������¼ ����M%��>�}~P'�bO~�,@%
&ކ�5���<	�%�V��{�qB)��q:��`����������
t���*R�������Cg~�)�1���μ�BB��u�D��f2S�^�9�>� ���#ӃG����r�ǁ6в�}y	XW���k�Z�~+�桑d"Q���J�Ȁ�6��[�Ҙ]���2��I��i�s-g5�^ؔ�I$�x�%�z��17����#"�B��R�L[�:�	e��Q�r3ӏ0X&�	�����u5�!�;���y.��9r��
J/Q�AD�})Z��=MK{?�"��c��u�0av�ʠf|A>�!�`���*_�b�x��j����g!����Fg#��V�J�Wr@���0(7y���
0�j^�B	|�?/��N?��p�2�Z�(c���f��J�}��?��hU#�?�o?wO	:�)��ޘjWU�u4gʯ��ˈX����q�\YoM�rt���3����2�%�M�_���� YN	F��(i��5��	eO�jX�y�X�����_h��*�*m�8�� ��� �a^��m�	��}>�5��:�"�{�\t���}m�~a��h%��{�r ��$�S��:K%'YePI\8/���"HИ�C�i	d�������|�̟z�K���P
�����6�[VEM)�3�������Q욨}C�sAn\�20�$�gF�˶�����{��CDA���W����1��O���$UB�����+	~i[�at�����Z������Փ��-��>F9��>Z�\�F�Sx�$H��k��[�i;z��i��]`��NwOJ�,x��4�Ld��XQP��2A�o�z�]�,�D��m�\���c\հ"!�y����f|vqQή=�g{�u���
qg5���]}��6q�QJ6�$g��Η�Q�#�oͩ6!�K��)��\c>3.�>Y��K��ވ�/٥�����t���
�4V2�%�`|Wa����"��h+�7y�#��N���R4�O��;�a�>��,�����,���YD1Fj�M.��x�M���+
p�(j����Qc��)=8��c"%�{#& �T��esBZ���À�C
�G;pv	3��D�9�<�i���uv��rpw���n���`��]8��Q}T�v��{lM�K^����zU�Y./ώG�R]�+�9�S���}4|r,�!#z$�n��N���[/L�k}�~1"+
@�yڋ�����|�4�����Fcō���ܑ�$��Z��T��?���b��m�aQ.!|���� �(�Mz�<�D*�z�g/��#H�>J�^��T�`^F�`����C�N��Jܐq;�-ሑ��Z�3#��G=HRVG�_r��h~��ZuuZD�J��;xy� �
��o$&�"_�`ضʷv�'���β��s�Q�m� �;Ե�}$���c��y���|�U���^� +}�g�<K�&�?����]a�*��\C��~�;(=�:������'g�YM�~�K[�w/��C��<��Ⱥ_�>|��F�-Δ?�බ	��n3��?�=�Ήa	L}�b��WA�.7��O�2=��KA�Yrs�9G��w�g>0z���Ƌ���������T�͉H�p���+t�d1]���W��}W��Lk� ����Q�h#{f84G �_~~��*�C��O�Ъ�������룿5�f�m�#��ؕէ$d�j	�q}�9�����	�r���Y_X`�=�p�!��6j	�<䬇K�Fu���b�8-�
 :��&ڇf��K�ߵ��ut5y�I�G�-ZSd.��*
E��[�nAG!�o��sd��'R�3[(�d�9�����L�5�=5� �W灤u�?)-�oE��JS���~vE�]��C�p��b!��-0Y�5� t,�b�'��fc=Y�;tݥy�k$.`��������^���F"K��g���P�j�b-�	<̾�Ϩ�D���5�{"��4�T��9��.�Z�t���"������m�WDϬ�`�S#p +b(���L����y���@�=������9�-ݽ�8��8�h�_[c��W�bLQuw!Z�%�S$�B��pV��XC�RM�4�N���6����VZ� 3���4�&AȀ���Y���[�3��|�  �u��.�kPX)z��ҕ��N�|U���"�C�ʲO��.�<M��2o4�m�b���Ihu�)�#LE��͙[�%H���+=�f|�^�Z+��N4��G���M��:�8#����,y7�����iT�*b��2��]��7Bo0�xQ�Q$�9jqQ:�9�cS��9`��}P�Tv����x;a��b>T~��T��P����5�P���N��X�ЈQ��'�+yܒ[rqs��$�)=�X��I/��
��ߕ��M����&ڥ.S�����:}F-��<)������8�ꭅz? Rn���k��"ٱ��Q#�I_�ٵ�)�_�%#&h�WZ��ȭ�57/����2����S�6m�<4�
Y\��KM���W#1��E���xn$�&�l�;Rϩ����-I���
F�w��Bz���Lr)��g->"J�Q{���+�H/p.��-�|��Y	^���w|�� ����-G�c�|�#P�Rf3���TZ(����H�S����,f�p����R�&2��P;�v��`�w!UT�nV�@��f=�#�)?S\�ဏҿM����pn:�^A}�<))��vf=��lZ�)���BG�͛�P-5�w��g>�tWҽysL�An`��4Z]n*
_��}�ۨ��j1o*�q�*e��ᅿ#���<6�\&�#Z �h/8߃uN���,u��$3�ƾ���G~�dg،�(�$���SR���S�la-�C7ҘI�?-? ��8&���"�iz�wM��O]�X��A�Of�D�N&��׌�
��1z-�� �����{��] ���V��	���qŠ���3�\熂���2T���Ի���*9��w9���~\c�6G�.�76��Eg���w%��;�C/<��=�+ڇfm���=y����ӺB��!s���F����V�]������t"�[j3.�q�#6F�8z��
W>�T]��?T΋P�h]s�3&}u��p��=o�c�g-(,w�I�mb5�s�%�r�К��G���3�_�S<�m����L7_`�����eV�cw-�*��&9#����\���Ј.*=鳮�}57a�S��ǅl�b*ȃ ъ��,]N��־mv�i����Z�1V#=�?PP�`���㞗��o���c���T�ޝ�a9�pfO�z�tЎE穇�뵗���Vn[� ��TgIG�[��)M���^lI����1_�5Sh��ri��~��>	jُ�b��a��V��w�Ż�c��H�����/ҡc�\%��ْ��X�#�	�����������6�k��R��1t���_�������F
�{G�[�%y��Ai�p�-��|���T�>V��lG����7�l��b��ň�Z븼����ț���Zp4�t��o���~�AbޘJ&�9�A�R�0a�平�]����V�"*��7�F\h����F �'�J#)�����E�?����{�T�ٻ���F��X��a����B�>K��/1h_6O{�~�����KZ<pсoCh	C�Ux�	�*#2���Z��Q#b�9�B���I6�Ӳ��^�YcMh���KΖ6Z�v�gHLB
�����~+�A�:��e���q���+}h Nl'���Y�,C�E�!�����0�����5/����ӽZ�&�'�'#ta�M(l�"��ҍ��,�|�Ū1�������_}��	iټD��1�"M��Z�&����GH.c�Ź��K4���:�K�D�Z�^{+x,���ֈک1 �	ˑ$�g]���n��>�|��&>�*̈́U�<��C��)/�`I�J�~�]��9X����ѬK��-ƪ��Q�с_���d{�H���ܱ��U�A�Q�_�X"ۤ�K8> N���ICN��Ab�A�%��{��&�(ٶ�1��ڜ�*QMz ��	�Q�߁zw3l����7��<�*���A��骀vW>�<��ebF3L����9�3`���po���ML�=�O�W}64�����$��D#6�H<��i��E&k����_Y�j��i�� ����u�W�ج����PZE���Sv4�u�t����wTN �%!�y=۲���(��M�U���U���a�c)��%;>�*�~ަu�4���{��;��Au�>z�\az��)�ɕ�Cmw��� Y2��æ|k�{:�
{��尴*m]�?.!9�v>Ù��k��r�
p}�ϫ���k���}j�,7�BȞi_N��/°xF�E�ăQ�BY6$��%��]�Z#�䦡�,�2dX�łz~I��U?%���/�D7E�8�HYRO`Y�y��-n�N��n��X�u��#{)��6�~�=j�;oR�a�]L�0�� zKj��404���G��Ivӯ��'.��:T��q{nFU�s2C�Fq]1�`S�t4/ZG����{*�O�ʘ5�j��x�:�^N�W䊛p��3?U5�偭�/�g{��7g:ep�{R�i���q2���z��fj���f���q�Q��A��n�Ne��P����9�ǀ����EӴPPM-\�F'%$ӵZ&�����i����=`#䚹���G�$�)�4�]��T�d���2/h���JQj�J�VT�h���qOO2���\~H�9���1k����X),z�݂�ق�WR�U�ީ�O�h�A^p�T�O�x��@���j�l�?��<]Π��@.�b��*��i�x��md]Bj�?�E]�B�>W�BL]�*�ޕfjZ�QđVP�nH�ΪK���- D��uX�@W���t��Zr� D���W���\�ݣ��y�YNp���Mv�󔢫�L�K�	��c�F�/|`���o�x�5�
���FLi1P�6���#ڪ�W���HӼ��!�<�ǌ���fp�)�����c��Ss ��qkq���TX��[0���yZ��s^h�+"7�?��������o��h������*�`�r���y�u#�U���C�<	�GC�E�9�>:�4o��Q^g���B0��i&:��*��~�$���Ih�j"�7��	1H� �:n�����M���b�ω7з3�Y@���?z����K�5͌զ݄Z �ޤ*[j��Jy.����-p
s#:�RϞvJ�
���t�'�(����K�ئL�S{2
z���`X����>�Y�y�x*3��n����D��j�3b�Գ��Z�t�l�L>3���W�� U��	ɖ��ź��M@Є�����k��b��X#Q��#x��a��\q�^�������NylKZ�8�z^C����y2�p״���"��f-�7�R9O��H���K���1u�)."=��9;�A7��Z
��1�v��yn{�0[�#}3Yݖ���U��\�;U�N��O��4V#�L����f��D��x��+�U�<W������-�k>K%BK�C���C�l,�`uJ�2��h �I:�/�2�fa�:mUM{�&���;�~ˍ�d��-���X���F�����
�G�$�y+MV�rPO�p����Uh�'�S�n�'o��c���/ŭSg���|6KvO��`c��,�u>Ϲ�V��Z�F�Zjǲ��N����w�~�h���![v�%�C=��ڂL�6|�̺�1$(�6R�&,����Q��2lq�u���3�yR�ٲ����GlIF]�ǜ�6�.P��������;���^�I8y·ʦD�%������ę�y�{�m|ȩu�*#6����l�W��qI�SH��6�bLG�a0D#D����J3����^LUp�	������@�4y�v��QD�p|�R��,�W;Zި��"�Bw�6$���1UZ�#�j0|ă;c��#���y���6qzNF��ΗA�"��[����J��yţ	���J�
��D�(���L��j�8MY�I�
�&n>��
/b�آa�g�����`���B}�tDB��+�?nwT����>������oW�Ҕ�ɶ����'�&�jgG�d��Xr<;��)���#gu^�x�K-3��Wr6�t�>��tp�r[)�놼%. ��PF�M�ao]l6���|��D�Y�����%y5��F�z=��+=�\4pd��a:�᫰Ki�yr&Qv=��5&���RO��8�MA&a�3�7i�5b]
�7�&>��q��7�P?L��/ N��B~�[3�GD��(�#f����hW�]�$��wF
�^&��żq�H`~3G�YQ���(c���w��i��5T���0q5MG�'Ý����q"_�$M`����G�3+{�N�<<)��7\�k�]�x��&�=O��5�:�t�ě�}a;�D+h^`��[�:�l�ad���åG���g��}�TD��3O�6�$�۝�4���4�.�_��	
Ö��������R\����O$$U*
�?�uA_(��|��n$������,N�XU�&K�YX� �]��.-���_����I���j���w�kT��f������^�ρ��[p�������$�|��NJ7�aRC R�H��<g�qv�(){fu!k)g�p{�W��K$$"��H+���0��E��sV���������ի�kO�#T���iyf��ex�t�ES���D��R�0V��rm���N���r���+�lM��y֌� b���$P+2���>8D :�hǯ��u�捿�ժN�#k\#�T��į�:�eK3�8��9�F�5-���e� ��4�2G�s��=��j�%��7�}	�y&MQG�o�4�
vJo���hweh�G�oMcd���#���IW��WQ�C�b�V1f��+r���C��g������9\fi�@w��W�%�) �4��2�kf��*ERQ�e�Av�8���9�����6�J�*;�I��7&�&�:�oVc�r䀣�w���>���g� n�y�1�5��4`8��$�$�3��*��a�����BqsB+2a�ʨ��"�\��f�!�G��>z�_Lh��y�vw�#��Zv�N�j�-4W�]'�����5n䥞�Y�xKv"�\S��(tN"e�Q��Nʉ�/� Z��F�������M8�O�]=r5Pg�z��t%�� a��󷼾���w���@�˵�y[`e�ߠ���MG�aybzJ���<.��%��h<�P�*dp�Aۨ�nM>�꫉R_�(�lZpM�WU�ěw��e�/�Hs!�{0�C�Gݗ_�r���ܼh���bc< z��6��"v�EC���W���!�;����$�Q%�^?�J��Au�cOt@�k6�}sO:�)�N$GC
j�(W�,�a���41yݳ �5������s%@u�/1�v!�_�%�m��>�{�"j��k	�H*o-�Z��0�h^��ˣ~�������03�?�G4�P��mM��,=�gZ-  �Ͻ4��£mc߾�C�脬�,�d����h��eք�Ly���/{����T�3,�����} u<R`L-��k����xq�|j��� 꼂�΀1��|��~$P)���Z�X�"�t02��M7GD�m�7տٴC��2�{����$�;��f�����3	�@�ӹa�q�/�~C��|z� �_�:/�d��p)KVG�S�iϐ��b/7��q��몣0��K���M�YF���gk����q|1��D�i����>�N:�8�Pn�PU�����	�j����������g�J�y��l�fʗ�sJ-M�hCj��G���U� ��?%�1aE^P�����9��<4Щ���+�dM�NB��C�qN�)5����O����m�R������fIg	�[�m�s�W�	-�2�q��|������^����1���8������{e�D��ȇ]�u����v��gkk�Q@Z�l)��D��3�YUb��b��~�"e�
o�l
�t���Udl�Ƞ��	�)���'�rA���Ye+�͜g��XՂ��'c��� �ۻ_���q�?��#:ѯ�Iv$�?�S<w�L���TI�+KmX�G�VLd=����X]��U�F�G뇑@��ҡG��J
P0n�[2
�0C
�s���<[93�pF���b�L�.���]����X䧓�V�V;�5 Z����4�u.�Z���ei����z���QP��:c_�s��d�tB�B=`<?#xChLU�`~KK�U�bZ��3ݷv�]K�jU�P���r�)��Ns�yT��Q�)���h�ǧ�Zxm��p7���i�(����w譀8� Γ����s��q��]�W�¦ˊ&��-"��6�	��r�"*��5o���BҁPX#��M��$ˬK.��?�B��R�[Ѽf����������``6A�����1{��G;�F�/N�z�H��Ho�jaj���l6�-3�ܕ��+3�LS���b�*��m�?��n��H���kJ�p3�?[;��x�e���a�j�!t
�:q�6�"��&�/�b� �X�2�|-�}�j����$�������V*?���k<f�k�GZ�"U��K����ށc�A:�1C��GcM�ޭ�$�=�f�z��oj	�L��dǉd��Y00k����J�v(�����M����=a�鎗A^���d.mkj�K��.�2�;(�J��Ԩ�0j|�S�B����3J2�eG�x�.�����T7Rl�z�^-ӏ���)5�����ʖc�t�^��s+t���F<B��S?�O��m]�زW���^
.�h�c�"߱WbB�ͽ�c���2G5����^�-��B)�s���j��!;ʰ�-�0����;� D
Cj��:GPtIrDd��ܑ=�����3�J�Äν	�%�"׋ӧ5�21�k����WY�U�Ϲ��*��z%w��d?�g���s�D�S�S�2�/��lY�F,3�U
;$�1���9 _2ɪ�����!S8^G@�q�	�������:d�ߌ��q�!�[���c�����)ro����5�Reo��G�E��E����OVQ��%Lk�s6KA@'p�K�6gU( [/v�4�I�fL��S�м�"��8��r���A���@K���}��f�Y�*s�$w�l�W�:���b��W���o�"��=c-��`��eS�M�E��H���o*���<-����}}�ΰ��5 ;?_��h#�`���u�+�� �S+�㮳$h\ߓ\?��4~.%����*/�+ؽc���n]D����tb�������fm�o:��;��U�,NvX����`p�����p�V<�/�-�&��+�K�t����c
#�R��+-S�]�\��}��HUV��X�B� ������>�W�� �>ӃH!s{zV�ყ0�x ���S�e����9J��aڴ+���9�Mfo^٩�9{z�+�~�~�DQ���:��G�,A�L��?E�����d҆���O�C]�G�g�4w�3��7������b� ���f=[-�z� XVM�i���!<goPU[1l �s9���|�6�wz�FȕN_��9��4;�n���\~S��z�$Z�}��+'���h	~���h�>�V'F�p}���Ig���+N�_�����Q �VPj �?l׉�M�m�b��C
���O'�!����_�6F��k����bSp�m�*� �l�ۯ�s��\��3���E����A�=��$t;/Ţ p���FQ�k�5���f�؃��9��aue��]:s�;]��/G�m��)J�������כ�����Z8����C�����O�� WY)k�6z��E��|���|�A�0���\����L+�޼�Z
d+T��YO Ay����e=Y�I\�Q��Kpw��eI̝�P��$���@�����q�=���Mk�����Y�����F"��/�����8j�.��@�6��$�!x[��$�r��+�l���5JE�\4�b�,���p�u�g���T��N|l�ʚ�u��%?3��U=��PI�{�j5�ct�S�wL.�͑���knh�q��?:1��*5e��T�J{�aþq��1�,*��h;�%� j��# W�X򦣏����������%�<q�ю�ר[�M�4�$f���;�zҳ}�]n��)�%[d����&��Xya�3��Ǒ,��5�PZ	���Ie�p���
yԌ�0��tqbch��B����vNs��[���HM�B�־�xB�(��Ei;S`�h3���V l<�MS�*�H�ʆ�O�n:�S^O L�)l��>P�{u��ܲ���e�K�L!�*�P�S�鼾X���L���p4տ��ʻ@�T&�dh��p�����i�����N@�Ez˒k��y�M"OD(��s�l��HQ������!l�E�f�6"Xw������j��P��P���΢}_\>RL�>p������"�������D����ԕ�A1黐f���D`��V/�u�Pw5�V�NƐ�mZ�����V��|��WH�p����!M4�O9�D���E�]#�� [�9��Q��96
�j�q9���>,>�������A2�z ~���C�@'�Хͭt�Դ�E��%�hh1��|̤�w�C�pi)�;m5z�B��}~�}���`�K������x�31���l|�ˮp�Xd� 6ݞ�m ����mւ�4��=��/���T����ړ#�;��.�)�g5R��.p7oY_��Py*�/�5�g�+F����eD���+��7cR�L����7��!NU-qŎlߊS	�
B���ڋ��g8$��� 7b����XS7H�x �>���:4jO,����(�(c$%�@!Ϳ�G��-�_bj2�A����W����y�E.X.|y-�����
ı$w�� �x�=�~Q0�k<�܄�R���Q�>�\�q��g5�V�	�l�݈ʫo�ɮ�5w����u$��tw�[�AQ�qܢ���zY�lQ6{e�w�z7�-�����7�������c�:ޡMRkL��A@��M;He>�����JP4��ƣ������x�7�{ٚ�*��2�nt�_4q�¤��Oުȫ�MQdD���v��Db��j�J��.�Y�,s���?_V��;�!zQ��v��2O����^�o�0o�����ώ�� aEzu#tb��F$���C>A��F��s盳*e�v�/m��G��A�}Z�Xv�-�wHE 4�f�LK�����F3���~�l^��#}�����P`*?"��ϋ3��w�L�k�=��YT,�����t�E� �ة�m�$�7��ying+ͤUXn�e�-]L����DCԄ0�c�=���Uh0fk� �����(�#_��,�i�g�΂L|g;D���P�V�)3��s����Ԕ�Y(��5�&ɗ�sH�Zz��q��)r���ʒ���t2����2�<U��&"V=FCB`�8�n��:�� ���7P��j��}2��U�8�}v/d9���D�{8��*�ٗ�([9Ţ��2b'��d�z��
� Re76xz� s.N�@����ac~� ���a���]`�Spb�uZ� ��p�lk���x[+�.��q���yOȚhpZ��z9R�������=Ն���x�S~��q,���v)`0����&��p%$�X���4��CP����ȍ�*�2��<�����Ǻ�:64����?��QUC�Q&9��m9�3����A6#�����R�"���G�\��^R_��r�b��y��b�`�E���j�g�Q&�g2 	�{9��@��[kc�}���HN�Z{+a飯>Fw��:����u(��B�6
�n�wv��2;�,O-7�e�
�ƶJ>%����|�~L���Ĺ����p�ǾQ�)��:�ͥY<�|�6�Un�T�a����i�wku���w$��Eg���ɸ�<�����^8_����JM�`o��:K�0S�D��zk*����۸d�l����)���|�}"�ܟ�ll>��-����W�d�7��34~Ga9ɛ�J��8��:W��1!N�ì�7]��#o�� ���$�#����O�h-������6�0[�CT�o����b��%�OqW-�6�V���:����q]1��7b!MXmH8E�W:+�m�����J��Kf39�'��d��d�`׌.r��\I&+?yE��onqrY&��=7� ��/ZRG=���*�->pe�.4٩�����n�t�i���x,g��쁽�"jDʗW����d$��DG���n��j>$��}L��`����J�d=="��	vt��W�	����,���ʦ0QpI Q'�(��瑔�Wh���Jh�E�����LB/%����"�[<�`C�h^����5�]�JIEx,��8�u��4^%����`}e%�)S���I~���������T+�����K��_��wN�<�_7�n&J�$c�YuZ��Uݦ�z�޸u��Q"��0��FR�o[��.0�e���@�p!2@�2y��:�(�<`�0!=Y?�%=W	Qh�S;A]^���7���aqD�*M����m���v�Kx[�>J�`s��v�t��"�hF[��t@E7�����v-l 30g���Y��'�e��מHEŌ��	��	��~�3�YN,o�}��Q�".		�9������ӱQV������0�i�-V�@�R'��c�H@E��Ln/�)jo����7���kZ��j��=d�/��
g����8k��8L`H4�=�Y���N:ph�s�k�s�j�c����z���Ԫ��>�>!�ư�N�G��8����d���ܺ�ͫ�/�R��z��z@[�nU·�{���Bhr�t������fs�&{z�7�&Z_Ʒ�d��I
^�~fl��N&W����g�v�TȒ�R2���֤f�y" �j�Ь�:���\l��%j�V��ں�y��"o+9AB=��Z���`�j�O���:�l�s��m�p� b|�� N�~�{�
� ��ge�6K㭕R��,��G���
��7m��'+�����þ��`�r�OV�~Q]G���m�����8�� V�� %q���>e�J6��{:�<�f��P�T��ȸ���;#�]�)@�p�OL��Z(bC/����/���"D��$��}�?��a�[�A�.8�9���Ӳ�|*��Ѕ̼#���FڶvBz��Va;	deq!{������$o.C�΁!=P�2W^'���׷���7��@�s��M: ��E¦LG�vҤ���KpB�̏騻@�d�R}X�b:� ���~ܖ3�D��������	l��E���ܰ��3��-�n�:7��[޳��P�,WG��r��EB���$�Pٌ��Q���N��.Ĕ9^[��ߦz���=䢽6�:��<5ꑏ�w�+���#��5e�/���6m��\߷��IF���f/L0a�#$�Z�ۏ�K����
���6�D>ֳ��= �,n�D���8�<�r~{����ϒ4�R;ū00�(9��'�k�E�4��������yF�����5;�iV�Ȓrpj�S�ԅ���O��Z5��e���yG)�%�� �[���/\�ֹ[X��X�s���D��C3^��H�<�*��+�&���5N u|�ҿ#�na="Xщ���jR��p>I�մ3�u7Yn��'�KCT	dT5��i��d���[�N@"���	�٤�0p��#���������Ej���'��'C��$��,�p9�pKI7����L�2*�h���~�6������u�O�b&�c�l�W^5����g�V������4R����);Bt�[1���*���%����v�2B��Ϥ�>��h��@�C�hX�P�4�
}'�։�Gk���>��q��JC�~WC���Uw�Bx
m������aӡ��G�U,��������LHs	�T��(�����M�	�.ugH�B4iBDK�S����Hu|`���)���cm��?�!��N����OU�u���h�=�X7P�q�D�ge�g}x�1��@���U<�9J��έ���g�-���iܲ�l�ں1m��qs_	5���T�g��M�Yߡ���l��t��Y���,T�\��y�叢J��`┽\W,N�o�}3n�=����^�"@�gZ�����c���d�$2k��z�����R�O�9;=[���*�`-��gTRʼ{f��N��2�����ŝgn%2V�ԉX����<\���;�+7����FˁL.�
WN�yk*T�`�WqD��J��#�f���T�3ΰ�k����P"k����X� ̤��E�*#h,��Vg��a��}l����"�w���z�� �kQ!�O	���c��E�,�d��C)1:1��Қ�M��up���S��K&�����c�C���N������ݞQd�iɰ��X3��H���i
�ϭ��_�[�
�{DGB|q��{�����~�aב)��:���="`Wv�8X���%@��7M36{�t����~n�!m"���m�+𝑻5Ј)�r[M6g�x��O���-��G&��O/���bRw�G��EtL����}.��~e�u+f�j�П��WK�߼��B����ܱ©���h�������.�����m4�$԰���{9�U2��C�D��k��j�v�{�g#n&��ԛ�����~'���9+�C`6�Vj�ͭ�*�I��r3^�ߒB�u��W ���oa����
����� ��t�{���⋼Qk\�?�G]t"N5T����B�	QM��G�����y�#ڡ����2�X?W�&�3�'3�"*Y�e�# �9$����b�A�}s�q<m�*���c�E� ��׺����3�L�hή���|��1���&��ʡ�2vĊ��`i���ڋ��I�h1�%�ςݫQ�v���$��N5�Jy&�D��>͍��|WE����9�xH$��s��)����нKr�9��@�mE%X/*���c�}yE����#g��oS�m�+�����o��ŝc͛�����_��r����w�RAI�V����(�E�9�Q��j�����b�͒�-)T�0\��L������O~�2�e]�s�
��!�y����x�%�8/��`�.��s�m'��&���I%V�*�Lh	�~�l܆�2=E|��݈-�d5����KD� h�f:�>���cձ˽]/f&$,�N����5o׮��Q�����W/�M=N"��9f	��MY}i'��"�Sg�Bb'^ H�)T��.�M�⧥��i�.�{��Y\2����=�����t��{S���"V��Ǹ;6Y�I�r�8�*){,c��x9ᲄ��1�1I�^�@������n��u���W7ف��j�,Bv{��-F�i�ā�*��^���+.wt�F�����LA|�R��S���Hr�rY�HB��3w��O�eR�v����Ӿ���v���qd���c(�	�+�@�}n�GK�f��@��\B���9����Dm8Ѐq��h�cҹm��Xs1Q�����5Q����?�����D�Z4|pg�	Dl'���wܼ
�xG�������B�����"&
��hH|�*k�g��avPz���/�/e[�X�x{0���aʫ9��QI]��b��E��j�E(5ׁAJ:{O&'���bƜM�9am�0��J�-�x��\��_�4{C����I�tn���5_�b���r�3��_
�m�ٞOu�c�i�}�`����%ؿ���V��e�\�a*�i�=�-̯�)��Ҟ{�a��i��i>�Tl�z�/�\n���H��	|��lz*Z�@�����kU�\�L�O���P ���P�S����?2����t殖%���Ϧ�AِLM�,�^֌�*�c�Sa����J��P�a�Վ�C�{]�CSY��3�V�)STL[���?���&u����t���a�,2��r�t�Q�[��ʆ��������{%G\غ�`	�ǵW[5z�J'��,�۴u��8j���QxE�]�]�·� o�2��薔8��r�n�/d��,�%Ì�g��A�W��e��!B�T����v�Ok��;[����D��5�NC�
����Cꮳ3��`��i�~WV/\��]ӑ\�R��Q���M[����<9௃Yq�q��Q*�k�<��$@tY��qY�Jk�=W�*���=���FӍ��/�����
�[۩�La2 �i9���;��~T��e����t#�}������M�7������4kį�"�����1@��[P"%V�i%~2��npr薓�{��5#0��E���H��^p�x�z� �m�%`3�v��&��7^�%"�J����U}0�(1�s���X��@OE�#�ݔ��r����G�Ȏƀ1��hK#f��&7~L��l�����^ZK��YdX��;l�G���!�U�$qnffs9&2�E��P7�g �hY����a�G�����/ٿ6����q�w��2x/*�9&"�\�](�x��Vxw)4	���Nl�_5n�r/>	O�� �����R�5+�.<�А�PHB�I�Qm���"?�~L���{����8��=<99�>;�ҭ��b�������?5р|�I�sd�F���*�1��H�Czz�F�|�-c�S�s84ɼ�ϡ���d@���ڳ@0��M�8�ix�!�����^*VH��2>�UB�9����~�YX�#<  ݄�W�iꝕZR���!�f���� ����*�TIѹ�����V�ݡ�͛D��k�Pg���I��($w)�ُ�	�����N`ㆿ��(�%���~L_��!�>"��(9	xqi^(Ys�tV���Z44��4�@)��uiU����h�(�(<"��w�j �["\K�(3uwĤ��)�g�ݕ��[��y������]!�]f����^����jH�֯��*�^��<U��Nd��@������ 0����=&i�rG�㴖A����� n��u���t⭎�&�5�?����%'m┟�0Z8Ce�`�zT���SVf�]��k�NHH��e���	,{�_�8h^6�t(�v��۰��w�s�b�:d jk}KG����:�Pk�6fE,Z�^������p����F2l��ɹyi������yIdl���8�lU��9��O����k_���_1;��xt.Vŏ�j�%�����s�	���?�Hpa0P��#���i�B��}�YoE/��B��:��3:�p�q���Q0�b��o�"i_[L������.��P����၃_�,5��LYq��+�S�T��ș�%�A}Ċ"�\�����&���kfl�WF���-�d�5����ؔ�a^���(� � �����+/��MV���~_�Ȓ`<�F��qz��U�T����[�#iM��ؘ�W��X���ҀTaf�;vK)#1����g�j����V- ���>��P\�խ���W��K9�V�x'�Ό\�U��$�\
�7ƌR���0�I|�jmW`�:�^����z��X��v/�U��(�_ڬ�:��"I1ꣿ/��v�
��E[��(4?��4kp��v���#rX0���Ȥ�F�h,�u��T��G`�^��ܲ�D����W�@}���Fg�=2�.^�ßFƉ�rvӘo����
��`ys��6�[;Ebt=�kE��,6 ���0���o��'���|.���:nWO|���:�����:ͻ^M�2;�_n�������;��!��_/�>��k��sR�U-IK�#?1b�Cf��4Aм�k�pA��|�x;4)V�����f������:�3�0�t�S�{7!����'�G8p��EL)����K��C3�^C�s8��Q޹�*ߺnp���/�����5f"o�#8A��>�*2�O;�J��"[J����F1����qi�$ %�nr�w>�-���tS�[�^VSBi��.?�Ieݕ����(+0{Сy�rG�%��8'Ҭr��ƙSFr��+-�*��;m��jǮ=wX���������Tb��;���|m{ tw\���Z�����e\O=�
Mw �T�88|v8xi�!��!���k 	95'ж��eb�F\��
���_��Yo*A^����sZXGD~HE�!�6����GP�w�
�8"���ɘh"����������k}X�#��Gc�td︻�&�R���0��b��A�; ���ux�̚�a�:������en�[\�a5����r?󣿲U�.�k�Q:b	ޔ{�n��p3uaN^n�
�3HZњ�������-�R���@@�bm����+�_��ܝk��MGƼ�)��{�Nߨ�"���	RD���h��ߑ�q\3a��T��h"(��
�v�zxr���&c�n> �	��~�D�y�/��ѧ_�G��l�$��Q���S�`��X���6׏~����3D���R
��*_���C�Y���l�����s�?��ۙ����U��}�*-0�\�bp�Q���sB�=�F>Q��Bx��,x�=G�m���QJS���/#��MˏZH/1g10���z��ܰ� �%����LlS��V����FI��&	��@��@����uZ2h��k����U���P�=�,�~h���|G\d��%�!*�'\p��49V� �N��q�-`�'�S��i����*$���e��]WN�����jGh��F�r�| �;��S������=m���^-��D��y�	�d���CK=r)�5k�}aF���I��td����bK�������"@m�v3����5��t�bq���%�2)�yG��m�d�O�a2���|u���d2�d�@@���N��È�����s��ҥ��L�`:p`+<�17� �s�$P�d�52)�|�l�؉=	�j6XG�:���1F���.Ypꮗ,!6r��<q|�՛����e
�z
������I(�Ջ@"�����9�O��-�T�|��'��&գJ���Y�J����*@Q�?&��PA�e�>�O �3������h�'^��qE�\��ǃ���${�8q�
�j8#ps���$��Kc�y+�l����Ǩ��
K��U�9W{����p^;����b6�J���*o�<7��_���W�ö��8)SQ)�x^fxxUoNYv�UA+g�VDY2b�op�Q�^JxW������5e����P�� "D�!�>EXF��=�>U��ee��}Q�LH�kW��P�Kd�uV;��O���u��	�5�H^D3����W~�l$'�}+�|�੽�y.�`�uw����@P22�I7�zK�֨�ƪ��?��]�.�g��]�TE������ �{��ѹ�xS`�ߚY(��;Y�f
5�[��6O���'���S�{���|3�6����	Ye���A�T���'�P\��xy O&ߥ�hC	����i���njw��¹��jx/�2ɶ�R9����-����/-�m���
d5w�}FF�	�$�Zi��ʯ�ڏ�>�a��b����1AH�$Oe�z���4��i�U���eTe&dB�ԓ�����`�OQ��%s[�p��ίT�(/��V�"?xo�w��g�R�P�W;�� �/=N�\��(_��.�¿}�/���2��xO|81=.�X���,@O\D�2.���; ˾A<���^�U[x�͸�\�0����bT��NM��+����Ú��*2�㖨�]:	)�-�d�j�����U&k�H3��Ԕ2JqG�B��N<��b�����k ��)�Z_QH��Ϣx�du�������ْ��')��J����Vԭ^L��||�prB��^D*L���?`e���h
�7��7Rw[��e�m���9��-�e���=Ij��]MzS�G����A&��i3��	�����:�cg@\Dk2�F���� ���%28���;�U���Jk휦�FR���D�em�B�q��4�"�4@����cS��]�`��$�XR�6�,����I<_A��E@�̘�ȢT	]\�¤�T~���N쭺��x��9̌f3M\E1ٶ빎�#@��*a�9�h��q��5�Ɍ�O�n[�cJLy¹���`�9��J�\*z��|�r���%�BDߥ���i�$	(�B�#phe8�g���&5�
��2��\�.7.�(𕢹j�
�~��;V�k���k��$�C'�����Rƨ��q���u��5�P!'�t��Ю[w�K�?�PQv��F����[��d|Z&�ńts /W<Xd��OW]���Y�Ē3�KU�͔/�v�r��?n�h\�|؁���g���񹃐����X�I�,�)�`����u���%G�p�L�r�%�?}��-(�7��G��r~�ve�B�� ��x���4�y5@7�(�(`]T���&Q�Hl� a��F֗��SB�k��Rt�9&�~�G����3��xE��p��T'���Z����%<��fՑ1׶�"E��oGE2�!��O�>3���o�7����Rw�^��r|�w�gz���S��MP�Q��+b��ɳS((�=}({Q'�1%$Ri� W��n���^����v��%����#r�,0�/(,��f_�ˀq�Ɨ&k��o��{�J��h��f�60c�~!��ob�9�Җ�Z�m�ev�b9q�cι
z���z.����Lh<\�E�����{f��]��	g�k��{���Mv7P;��u3Ӭ_<�q���tn9�� ��� �(
\U�%iu�X	4�Nm`(�
K���`�H���??j{�N*�%�7D3�����(�e�9 �X�xe��z_�n���\�,�LĎ!|bɔ�)y�����'�=�Q8�<#o��FR�=)ջ��"z7*�F��˭Ѓ"Q{-B"�h��E'�+�]3�����q/g�<�E�p::���\i)�;���zl�]��\�Z��b�1��pسl��ŘƼs��� _	���N�˙ ��F^h �n�仏���T
�,.u�	�и�C�m�1@�5Y�ĥ��t;4m�3� �W�tT��m��g�x�V�c?�ߨ0�0ںxy���H�������)qw����~�~! ��=g�g2��!ʃ�+`�D�s��* �}a�t1(�h]c)ہ����B|*u'�I&�yc�������T�w����R(5��l{�v�� y��W�W'�3�*0A3�ڨ�8����h��Y����[1 c��hn�B��C�xw��ɿ��k��׻����kͤĳĿ��J�8&��OX��E\;:�
��C��/��q	p�|h�=;n���q�%t^�s�\��]'��C��_����FC�o���$	 8�>H�`�g��=;��셍�m��4��߬�8����o�P�;	���7-��!�KJ�wKd�zj�>7��eܑ!+���#��:�&Š|�!Qr��Q\�J!����G�qs)��L������a=�d'�wd_u6�Nk 0w�g��v)��e���JH��3(LǒieD�Y}o͈���7sy�vN*��Y���8@>��/tx�e���jm���׼+��іS��\�ʄm���Yy\�T�1��Z�:��Vؼ�������k&q0�K2�`�e�4�՛�g��Im�Mr�C:��y�cz���t��q���7>��(=�Q�Wy�|nLѸY���w��@_B���n|.��ú"`U���5�vS�e��0���Ř�9X���.2���EsC*����C�oH}�ʢ"�!9��r�p�9���j=�`�#����!@���*(�	A6;�Y�y�Ŭ��AR��Dvȑ@����ة�TI%��՘*G�Nxn����ՙB�l#�|�UcܲF��2'�a����,������&��5���4�u�l�P��fj?:����p?X�wY�G�L�;W6)��YZљ*Z�� ��r�b��l����/M�Jg&��FɽH&�8���3c�����M��"#}�%���}~K�A�Kѐ��>{����N���ZA-弬�Ԗ�kQv��9\���Z<�#��P"�Sp�ЋސצiقDE"~�۹�,�\lJ���a��AT9��n�B
�+(A-0�`�n�T{��Zsv qsa�����"�{
y:w&�t��u�~*bIח��r���#H��W��>Pu�]v��X:���;)Ey[�?�8��1�e��x��u�u��ٟߕ �1�ғ����[�㢢�҃f�6��^�d��(�z�W���`�)�,�H5��Y��	Dڛ�S�(\e�����2�OQ���*}AY
T�c�p�V	��f�-�u�W�AX�ݺa��ES�!_����`��hV	���;ߺI�Tn�B퓵�u,�X�^�*j������Dz7��V,MC�Qa���x#.E.v.5k�OS;�����a7(�������(+?(�-j�̻!W��CQ��a%<�[\�v�FE���5F��B�-k'�@�.��ַr����� .�ua� �`�([�"í!���PU��mN��K��[�|~NY�ݟ�&�d�0ZkEս]��)�gI
��ioba亭��Q�ߪ�P�����XI�s���I�;�mZ���V��{���=��B�� �s}�z~ț]O)@�{��;�8U���m�����h��^��������}�յƐ��7�@G?�:8��j�jH�f�,��}��}�Q����y|@���sC���c�q|�\�}eX�M���dى2#_[@����1v�o�*��V����d��D�`�M�w��-�J�1�H�qAk��(R<	�"�-�����5����rS��qxyу��;��=�������=��i��y�n;vpCoz����U�Bb��tÆX8�T�����5n�p�����iᘮi����8Y9�iad�����:Wa��3
���,ԗ.�F#�<̤���L�0�,P?��ų�]�Bh������'0�[��,>���e	������t��w
4�J�Q���1Kl)x�H�_{n�~��cR�x�%Oɝx�Q��E�Dx�<��*��9���檍�=��dE�)n��L�u��uΎ��	�u�A����p9OC���m7��9b�D���DŝL	��oט2Uv�������� HX�g�N�4�A�NmƜ="N�c	�C\���F�K��mY���ti"<\�[�A�e��5
�3�v������{��xH�rS�'YS9mYPq턑����}�2��m�?ϲ�4��d1X�%�B}�h�W	s��G1/�3��~�>����#t�h��/�=���h���,����7J�Bta�9]������jѝ ��� �X�Mx�����#�J�F�
|g�T�X�PUf�o�6�'eJ��]ְ벾�>S8f����Y78��C��o� �M�gO��r�1��r�%��`m��}r����9S`��3�v���_߿O�BMT%}6t�Ӯݽv��G�T�la�U�2�ԃ��ݕ#��;������s�wx��)-�����p�͐�ݽ�H-dTɋ�a�Dd?��d�W�g.ԩo^PXBwI�.z��w��(̋8�.���,M�B!��d������o<�_[�Ӌ�e���S��-Lf9�a�zt�KLMW�a�!��MŅ��e�6�]�{����K:��Q,�gj|}ۙ~�l�#Ṳ��HX��oI2�-�1�y�"����M�R�:m'�Y�)�T�mJ�m)l����V�k6{^���b���w�:ccB�*����7�Fj7콼S6N�Y�i9rO� J�K��a�x3����=\��>��#��	^�L�� 9�Z`�w�74��9� �S>��yn	�W�(�<�nMQ���(iԉ��f��m~��څ��H���w0
�E��̃�
S1O�jf96�v� ��ӂ 5ynu�@��֫�{>?��xyI���Z��T?���g��m&�JF@��E�'}���o��x�:Ұ�?�yS��6����Fr$h'�L �&ѳ8T��4�7ֆ����DJKDw$/-7����ٽ�8����H*�ܞ�_3����"��hh	��M|���4�p���;�j�E]V�!ݨ��ժ5EɖD��U�K�W��Ǆ�k&�$U�zZw�| )fH�g	jol5B���99�RT5��lK�����~ S��J��,P�I��La�cW�5Nu�o7 ����'nӨK6�k����
�o_ތ��*�!|��)�m��-�}�R.��~���[�e����Vp�� ��c�F`��Z��[�إq�v�+V��1�/�'�C4i�j��j��v�/�z�yu���T�Z$����m�|o���o�<fy���a.0�365�z�ВFD������!�eF��=a7�,d���ySdO���ӧ��OӢC� ;P��AYt�#��'Lә3����{�D/�h3�D_��@� �;b�E��k�ᙹ�(�V �R�$�eF#�־��;n�ճY~��FYr��ؚ�JG 
�V��l���	�0k��j��>H���8�7�ޛ�`	���"b�����;~�$�3�`I�0�����/#�6��tZ���w0��6U��=R�*�G:]h�&Uf�n���n�'��y��w��U_4�`�EcL��S���ۂ�ѣ��;HP���9$z�!������	�}��P�G��m���8�}1ň޹�����}����(A��[\�d߫�i�*��[�1���.�e)�����VL���e��+5��A��ȝ��0�*İ��k�
w�$�^���F����b�Q�3��+X���H�vM(w�G��:�~�U3�㠜tt��W�l�ml��lyvH��<���a�.��-�❸���Yt���T�k��?i�}���إX�K錅M΀�d�N@�]�������ݑ�d��Iܪ)������Li��}�U�1u�RD`S�&N��z���
0������2���?�Xމ�ҡ�7;��̌�RB����D$�-��0d�>�H�K&�����q
����.2��R*�D~[�!ꆠ���tA	q��7�@�E�V)��su��՛xe�� ]��i+x>E���;�R�����ԏ�K&�ZH,ժʓ�I��x��}a�u]����U�*�i�ɲ�U/� D�s��J�j<E���X,l
��4(� �Gn��v�e}y$�*�,�l��ރ��x�$��ox��=oLϽPlC���1��~v���=��xUz��f�Z��ǜGx.�{�e+g�\&�O2b]F��7����`t�6Ql.ו:,l�vK�:9�
��uX�b�h�u�O��u�E) ��IX#�UdsI[&��w.K-���ݐ%C�+� S�*�A�" ƂS���V��Upޱ�n)�c�\�6�Z��#�Sᄃt�a_`�^�)�%�Cf�*��<���4#*\y1�����^�����!C�4x����V����E����4��~����q�l�k��aШE�)��z_����̦Z��`��(�_k�ݸ/�]�YpZo�P�(�w������攸�bʀߒ|� ^���0E�	5b�p�(19�"	��&
]�!�HU���RX�ϹS-"C�:�UW�d�C��}��ч�����et��w�]�Va*c�E�a�]]ܱl�i�T`ܺn�)P>F��g�U�8�g2�ȼ5�1j�l�A����˓�ܟ�f%������a���J)�)��(����2h�
�(�g��bx�Tp�k��8av������#�ov�8hb�e�aA�y ��Ξ4��W9�ΰ���TGG���|�v�Qv��xAO�kU�ڿ[��=�h9�;�<v!����Z��Yӟ�0�y)��9����Sw�=����H��`��.J8��Ҳ��mT�r�Z=}�@#)F����߫-�4�<�@x�c�����k�'�)�b���BB��hy$0�U7��F��,?6&���JH{PJ�����α�Ð����P�)p��q�� ~�s��c�W��L��ᑙZ����o8�o�ڧBs�9%3@�W㊺��G�*�m��xSlm1���x�,9D%����)5�R��)'��t�����G�E!��8�r뻰$[�>E��O:!i�����~Du�>?���S_p�V��:�_�É��K�Ƅ�XYَ�����q߰'��i�J�tTǺ�s��>�6����\���Q5 :M!�/���p�z��x�tm�(�G�k^.�t�z��*	��:yxRl+�Z
d?�����">���sD:����Q�Ye��f��B��Y�ɟ���pv-�0V������#�r����.Gt���3ot�Y����~D��^j�8��Y�|B���T �v�#��`��IL>�@i�{Fh��i�����.sT���9�:��k�*gN���vq#̻��6�r�ҽŘv���y���8T`8@���P��)�����њ��%q��) �O)�����4@�|A��7[��rOl$�ʦ�U�60	�8\�\�gO�]��0|=�MOQ��5���Bf�z��?���������S��ĵJq�o�gCߢ�`�n��B'4?�9�<�q��Wiv��g;,��+��nb��o�P�p#X1�1Z*���a��r���y<	�q�u(�~U�W��d(��K{J����x��f�rXF��"��������mX>,P|Q4V�eB���s���d�z�e���f4�.��L��Yx 1p�w�K���A�"�rPww� ׶\*�EG��.��k��878��d���o��y�Y="<6�u�,�����Q�24
NE���:���۠|�F T���pX)�iW��mKJ�XG��j7�[M�.�E��qZ��'�]��V���i{�rB�u��E�����^�|CF�ұ�NjD��0Mz�֯�Ml����
�#�\���'k��>t��<����H�8�ͽ��'Hf����!���~���h�C8"	 ҏ�޻H��>�r�
����޵��vDm�G[c<�*��:?>2NUP'h�A����`�򄶹���s�m5��I�������Ydq�Gzc�Ib9�Z�z@���2��锑�P	��	
!#	��������z��Cy�{��i[�5�}LK�����j���6�p~���}M; � u/����I�Y��[+�(7��&6��nI������\�B v���!z
�4�Cr�}���(��޵H�\`-D*е�	��2e��J&�(	�qm\�w�\p�c'?��D�����~�c/����"�0����.>gD�/|ؗ��{|��u	�J��F���,6�8�4�VL����=yD@��-b�o$KӮDu��4�I~p�$.��[)?�ۃK��6�/�s����M$��ހ�&����i�X95\`���s$⾾�	�j$a��&�J���7��*1�Rd�����^e��JLL��zu9HL����V(7d$55o��/��b[b�cA�
LD�Wց3p40�g�o���S���g��.��Sk�H�� y��qb,��vΙ����\���U
BAz�WȮQ��������_%(i@��C|^�����&
T�NC+:�f��`h��TQ�E���[/V���Ź�)�e��ᡄ��Z�\K���B䝏�֑-��Z��s�`��#"8i8r|�b���&r�O��C�U���_V��G;�m�	��٬�-�����쯶�-n�e{�2�r�~�伖~;ݲ�ʺD���x@q�&��Y�eXYu�_f��J�k���d��j�X��k�S�?�AZt��>��)|����r����OF�#ٴ�x�{���5���;�y;+\�\��^@�K�'@���7޹"O� ��֙є}�a�9�e�v;���`?�{�̺���8����EU�����1;)%e^��~�c�Y
�园��f @�g�@e���P�Q{o���*H���e���BĶ�SА:�:���0?�p�9{-��Ws5I��;1�]�^�Z����^��/�%�n�$����� Tk�f�r�S	W�B�1�� �G���5s��j����P���	3�)y��7p�'���C��'3������xX���=�PׇC�TH���!��Ft�/fn�w�R��Rp]d2�ΆV�5��|�昹�?@Z��3:���gn�m��8F��k=���wp_Vm� ؇��i�N��	6x	�{�&�����������wJ�����e�1ۅ��n*�֯b�M������W�f-������f�N>�b �&���.�+�V�ô���f�~��p3��FF(R�+H�( 1>cZ�(ݟMu� ��.tDLR&�$��p�R+�nї� ��Q��:���TֳM��+sn��3iEKÕ�;�:���Xԏa��9��͕c�p>h����Θ\dG}����f]����� _��q��M��Ub���=|&�uh}s_���#�Vě$Ӧ�dIY(Z_�d]ј0B�fi[D��A@Ю!b�n�џf�K�n�X5Ƅ�+���k�2EQI�S�<�<qe�}��{;��I��C$x�r&�mq Y����W4Ă��xQ$"��3�Ѥ�<q�ĨT�ړ6�Zſͻ��[~�{�*@16j/k�a�f�nGC�葑wk�r��M(ޗί��j2"���VV��>�z��:��-wy���ń��S+�{�XÕ���m�ny�����P-"uU�s�	�ܮp+�!ާ-n��uFN�/�%CShLg�c��q�05���t�uG�B�vY�/��VaG*�ҽ�J�d�`�'yÅ��Hd׌,xKl\������[~��)냧�k:����Nx���߆U�ׁNG t�Lۊ1����,Y2����a�c�	X���r�Y�6�ae�.^��hQ�6��߭����s8�J�ݾTq\M�l˵���SM�	7�ҁDv?��5r9��~��K7�mY�*4��
�0{�i�#��{밹ǭ�s���BTd��M^2���IǊ����19�!d���y?���_��,oҋ�N�{����zm�Ǘ# �/I`�hG?�m!��=<���A��4���w��P�iB]��*� w����.�R�k���C���1;����N���_��W�kw2�B$�5�6�1�!C����{���c�W�I zٙ���:t'��c������X%�;*��'[�
}�X,D���e`�mB��M�5q�� ^ݰ5�R����h�[�Y��Bb�u�n=�`��pQ	͞���t��!��4[>�C��;�\qY����������y���o���B��
��mR9�C[��A�E׻�y���+	���T�.�f�\��e"�O���y��r4쌿*�#�@�SY�����~y�?���r�b��������T{����H�a��	ٞ�7��o�1������`�3�|��@�p��!x�p�+�T�x�aɬ�֯�}����b+��w�ܗ�s�oQ���^�.#ݽ<�v��E��L{W��C�*�}|��-j��|c�u��c���N�uBz_�RN��J#7���&IV�D�x� L�'���Áta�v��s(6<VE$'�Z*I�M�3҄GZwݻ��z����C[:n�]�g"B���\Bl	�p�M�=H�50�4�
��2��Ω�p��c�����\�n��GCܜ���dH����A-�C3ٙ�Pr�$Դ<d3��/i�ʚ\�򇻎�PI��O$FT������6W�T5��M]4R|}�x
њ���(H�1��;��.��y�!����!�b����oi&�G��,��ԗ�@@�߫M"��qq/����x�HKo��f*f�8X��KE�k@��i�� �M�yE=,X�aZ�]�zZ���c4MhVp!R[z=��f`�#���Nh?��6#���_��м:͉�f[a�i���*"fo�e�"vo[Œ����nr�qV�����X�*��X �w��W{P)��Q���:nY��b.=���Qx�+
@S�p�Y�T����PO���Vѭ���A�+&O�b���ev�zn��5��:�@0��	��@��!\�0�K�� ���9�@������r��1v�%&=�])Jg~У9�Z{f�Mݧ �����70e���G2�p2Tӟd��0H<>)��GFU[�� ߝik^���z��󣴾Q-��p/��_7HJ��ɠP�m�XX������{Fd��|�
�8��
��q�\R��K
}�!�H�s����)#ּ����i��m9r�V�r�
���!sa�cw|�~��ø������9�Wo�����a���	�`�i�e��U��ĥdd�V�Ať���D���䭀J]�5r�,c.��,a|Z,K$��"���?!Z���9�`�Sީ�l�0ox�F/�^a-�̊�p�7p���^9*�gRQ5'܆vmr�F}*}����J�ù}�.h�*
���dX���4`��29�)�:�
���X��Rm�|�O��s���i�$����(ߏ�[��Z�&v�Ǿ�
��E.㴍2�ꅭ��<�-���\2sCB��ypf�������O��n���5 #^��Y@�5Y>�3��C{��3,�y>�H�p���;�q��=���zG�4H�N�鿬��ȓ0dq��]��P��,c���i��^"yc�['u[�ǣ�(�zY��uC��e�T�_���Υ]��n�/l��|�����X;�b�ۘ�C@pJ��E�li,Mj� Ń�x���&�+��HU<E�V>�_��J���%8U��_�W4�9]ԓa������Μm!Vs?/�i���������g����w`��A_HX�������E�M��BL��3V$����JG!(���2��;�0��K1:"�6�q�W��C���X:}_���kv�)6�����"�?��d���i�҃��9wE`h$aO��c5HG�H)�
 ��q��Ѐj@�J%s�mN� *�-?x:��L�Nz��{����8���z�P	�p$B܊BY9�v��4L���Ĥ�1pS���Au��u���3�#���M�&��s
a�θ7�n꯬�Z�y���6S���1�4ZH��r��6&V��ד��04t
m��C�j����i�����QO�ޘC�n0^P��� \�h�u_E�p�{Wo�u�vM��$�םL��:(�C�V5L�=F����T�d���.>��|�%�Vi��|L;��i�� �H(mH;Ī��{�]��,@�ષѕ���)`W��m�r�lӤ�y��s���{��NN������:��=��۬3�e?�b�Z��M[�)���D����YW�n3�E8�E��E�,Æ$׮q����G�۷^��K�%� ��Q2^i0' ���u ���(�`M�z� w~�"��P��9��fDi����6�����([���6'�9Y�H����n�q-��׍��ɮ*���@�;}���	�Øp߯���I;�v�m�	��˄�K��򮚁1�U��Mq���Rj"=W�]��Lý���8��HH)��G��pB��߄���9�
g�&1߸�Z&�y� �T���D���`ߔ�
G�!���ZD�+�ܖ������6"�TYt��>���$�gPvsJMa��0;R�&�pČ�w�B�5H$����C�R?���gᩁ
ƭ�"����]�7(ޅ�~R��a�Y�$f�E�EGSP�j\�+����[i{T�J6��>��x���e3�M��R���*�/ ��O����A'U�}tM #x��b�ۆ{���so�^QJ��P!�H��&}����8�s����t2��Yk�D��c��3�U/���8�����ΌC^��"��p�4��:K���l�i�����e@���N�4�|��c��}.jI�ɰ�\��(��~��N�l�w�bM(yG�[���9�ϧH<�QRӤ�D���O����)h�����C&��:c����w$���F0���&ú!�s䝠P��zFo�y/�xx�S��h�9]1 ���2�Q���o��d�ΐaZIHS�\�p���ԅ��`��������`����7 �ir~O	����S+�ϯ�1]��ɤQ�k¹LK�"�Y%��D#�>�Ʃ�@l�[�8��D9�J���-\��=�T�I��J^��RU2^:B5���3}Vne�'랶�X�Z,���P�2Z�We$��:�	u8�8I��wh���_N�lɛǣ]��[od��sv��?��K���B�IIN�[����Iʛ�[##[��+\@�C��V�<��ҥR��l�f\�;�mH5��5Kۢ>4��ba��ُ��uØ��`0�G�!}W��9R�l7�Ϥ�%�2�_������@X�͍�&�]�)�]�1����s��^b§<�rQ�y]�&0O�b�ubw�a�0��C��.��)u$��0˳���	f���g��k�.�����q�e��=�����ܽ({�����Oq�.���%/����2��5��\=����H������0��cqtl�vT�+��v��Ě?6���)�4�����Oc����	]h��s�/ӑ�(��hl��@Ii����X�*��%��䡂M�[����r�	�z��������g�Z��LR�~����>\�Ö�J}����&�q�D������48�b[��;�!�A�9��k�εt��6������L��s�2�Q?Z) /���Z?S_y���m�?��mޅZ�as�DM�B��C#U�e�!�L��7Ay�No���;|S6���:�0j��eA��k ��]S.�`��t"���`��6��t��K��w�A���o��ƌb�n^��	�i�@b�.@�pk#�\�D�����$4(򜟛�÷*ժ~M�0�?�qS���VW�pF���=(�\�����������ow/V���;~�[����)�<�C�Co��i� IDZ�p�}@r��xR�`��gҮr�A����C�C�Bj����o�Ϗf�o!P&R��1���%��YY	�Gu*~Q�8�иD�A��M�)8�Q�%��cS9�zˡ�7��K�e��}͌�C q
���2w8��/���¸ކr[{u�� ���}r���B�u���$=be��Dʷ����D�J��e3b6�9-l\AA���Z{+2�)�i�~wA*��z2�"|�"wm2�ƸX^�*o(�f[�)��l<�T�^�ÚH��$p�O㦱�O~-��ۯ��E�o��b�X���6v���!�0.�5�w�T�BL��PN��ER�,�h�^��M�XN������Vv��IJ�9��ly��p<9:n��3G|�'�L�ؼ��,��|���3�V>̲5E#�*�N����a|�GO��ma����֐,@Б5k��@��W^���v�� ��b8��R��E�n^�x��u�4�z����r�r��ొ��&󔅧���a����黋�C@�,�`��v�� ��̸óٲU�!*w��ߤ�m�X��:�~�/ս0��+��6e�������,v�����h���%g���og	|���r\����U����]J�Օ/fG|�<�B�=���u��(ǸM ���]�c_C���i��hN�$r$z�In�LF��&�����]Z�Y��^B���eֳ��AufV�{����I����M�����يQ���Hji��>�����m�\������ 9����dT�bB\�W��+���ǧ�^��.��}���<C�z�W�̹��~!
M8S,�ġ�!�vN�*��p�6����2o'uWq�V�iE�<zr+j	�g՜D	У��I)�c�己W�I�zƜd���"l�`�X����	""F����Li��\|�J������'iC��� �|�-=R>�PL�]Or3`�� m�ڣ���Ц@�N�A+_�cQ�unh�9�`V�K$͸�O�VT/�&�3Q�h����ͻ�v�y�W2�g��5�N��m��&�Q�&A�y��I�;EI6����i��
�ZQפ�Ӻ��[K�Ŋ��s�S�kݮ��fD�cg�58$|���{8���#��|<L�7'���M��x�W�[����Ӆ��(f�"�6X�~Q�8z�[|c.�%�l�D�����|h������L�r;���бf���S4YT��duYo
� �zDw�8����&_^KT�u;R�HU`�Z֟�=S)2��
��	:�uz�[��K)��8��@]������12�j��g���/�^*���cV"�ǼKr����A'Q�O�k
�C��:'d*�Ai�ݨ��;Rǿ @�jT��J�!�_�ՃVĂ#]FBy�t����ql;꿡��?�E4��k��y�| �9;E�/<ɼ��p��UM�������'5������Y�"֖�mrq������v� Djm�-�@��KW8{��9U���y\�y�P��{~O���+zw[�Xq����DQ��	�T��R��G����yk�YF;3µI��k~���J�c��O����!�/���o7�m@�;A������R
+�!��dZ��q�޷z/����]�,�5��$x9��:�ű���o��̥��i�c��őIr#ycKݽ^D�:^�u$��	��T��D�6FW��ۣ��;{�\�XcI�cDմ��7�DL�hQ��>:��3��PɎ��=�ʔf*dJ�
��I������2�rA��X���Y<��q�iY��yp��a����megy<ڤ���ڑF�4U7Q<���Y�bв���)\��fOM|�SΣ�ʣ��=Q�^��?_	�	�{���<���f�\0�PKvZP6Է�;�E�4�R�����6���؋=����%-�&�����8?w�{м(m����̏g������_Z��}�H�%=8W�����k���BUN�I���kH�������O?:�;I��#�h�"I£גt��]�<@\���*�7PO:�������kD��w�y�x⏙��( XM�`�B��#���1AB��B��(��f���(��d�vxۖ�3��ٵE�>�KW$t}��Ӕ��K��m~�]9,A䳎$|��}Ќ��[���drU�7��[WpC%~��
O�I"8�/�0����L�V�#I�"��E=��Urۃ��V�s�9���\��6Σ$���Uv�H}�R�<8�V�}be;0�l�e�E4k>J�Q�L��6��/f�i�(Tm0�Q-%�������� �6P/�ZLZj��f�������5e4O&���6��� �;�4��9�ԊiIKiD���_�BYG�G��CB;�Ђ֨�O6jJ�� ��S@���htI�Y�]_��%n3'��M����r�������o¡*���/_@���Q�
Z]���Q-�}&��&EWX�@��D�2�� ��..�^K�������o�U�wt(Z�f�-��(^
G���le=��V�셏7.N\L���;���+�'��Y�mZ�c��q��� �"���V�L9`�"�ǝ6��%��ڝ�.v�}㝓�<'��ۘϕ� ��/�2#��iye�
���o�\���ƼFRf�G�>S���ȧ�9��R2=0q�����АR|E���{Hʫ&j�n$I���9^���2F�����6�IjF�e��*]����~MI�Q��̾m~����^ p	�0У�N?�@�}�C�-��k�{
)S�3g:`�&n�bY�4�PЛ@^��Yv(��D:î���3���N^��7n�m�]�D��8~_2$�
�)�K��]%Y*��yl_m�WIJ������<��@=�驮�����D
Y�m�o�L�����]a9���$�
�G^��A�Z�ߗK��:��P�>�h'f�[�1x��U��h	H-2�W{�0q#��#���ͺ�} x$�ߍă�1R�B�/����B�r���6K�
�������@� Jd�XF��oV�v
rk3x�F'=���#):0���^�	��t�ͳn�DZ��iL�^�Ѓ:���-@t�65��/�����������Z66-)�u�1ac�թ��2ˉ/���'<};�J8������J�pT�շq�QV��DءeD&�83����wQEN�g�jW;��	mV;�IPd�a"�dv�n���v��k��塇�Cvt�zi	�D[�8�Hf�Lk��&�:h=�VW3����u�'�� 7�L�t�W�-�^;�s�.��}p�3%� u�|�����|�9\a����ࡕ(Ēy��\�[��(
13�V�N2<�$H�iaݡJ��3G�����������$.É}��}����p�p�6��Z����&����
��}G�v$c{8��\F�i?-��Cf, �+,0ؕ4��cE�+6-�C�$����?�N��:�4Gg�$	���&���Qcx����YE��ŖF�Q����E�:����F�>\7w���b�jb���It3����B�>� �Iv�EO��44X��􁕆��3�UI�r�h<67ʶ�L���4����t���ްb�H�n��k��u�~�FA~��|�O� �sY�]�i��qC;���P�)�
 S���48�%�]׮�Q����ױ��͸
�n�hٸ���$C�7SqBD����������>t!�Y���Z�uqd�����z_�{������)���j*��J�̾�����'NS��J�y���x���qR�P�!UТ<����4�q���O�'��5���; ]�8�>f_��}7T緜��n����6c#ZJ��A���F�@����׆O�z���=�a���V�U��x��e�0�+9t�b!�Kum,�FPEZy��i�I��QǊOP۷`�Mg���c9q\pP��`�x��L���'��N� �PC��;jrc��H�q"<A�MdU3�������4�h"�hm��J�q�Q�f����q�Ϻ��6Rh����?�"* �TBx�❘�b����U�t�����(��"�-��/� ��ۍ���+1��mU��~��tн6^:Y����4�,�m�=��ĺ$�u)�GP��Ǯ�#�QB�����q��g��� A霵Ŕ����;�����74I�C�j|��&�n*d���\'"wI���w���!�͘���ή��G/Ʊ?��	(n��y)H��Ss~��e{�&����@	�㤄���pkN�*�C��K	�/�B�1K��	���z��"j���u�_:�%٣�e��7�p����\�ex㎳����B�p����~ �n�)�Z���G������mp��z�*�g��_$7IR���pM`�&?/�lLo��N�H	Q���WI\i2%Kq
�P�|�^[tP���!���e\���k�5����T}]M$R�?^]DL�	�E�6d6a?�t}����`�iӧ��ED)�h�0�^Jb����䢭��uQ�WJ�w��9����-����CEW��i��G�[/t#ȲG��PQMmUṁM���@F�	F��l���=�A��C��1Щ�|��-�V�<k:�^��LEZ���Tt�k���p�B;�RC�I��Q�R��0Po��eAtw)�����S�e�L>4�t�� Y�H4p�`]��|�����;"3�Ф�����F8�w��>����;�a��6�O�`�q2U5�M����lzB�U��D(�*�����&�9�����IЯ2W����Tc�-����H�ԩ0gA4bG�����Y�o�ֲ��vJ���a�'R$�ـ>n�N����j��E�.􍷴�w����Ҕ��`�mZG��^�ۄ@=ҡa,�%�����A�͵�1_��H�,���@y"�=>�6JZQ�8,����l I���ugB/о��뮕�v��h��-_����	�m��,EMБ+�_�"����EבV7 Y^�,L*k��0[���j�y[J����5���0�M@�Wl䜡��1>}D�)��~&X�J��!��5���b��ɒ[3�DH	���n����L*|�f����r
�W*��L����t�M�O���r����s��t>�o�LJ\� 'q�biC'������1gg.�KI��͍*�@���Oc��#([�v���%#�u������f*��_r:�t(] _�
��U�n�Ľ���E�������<�v�ן���jo�&%YZ�`+{��>�dݏ��D:m�G-J��%�/�'��k",��UaS���v��e����r=��֞�j�zQ����K_cz	�a6^��\B	�|�+.�yQ}8�S$���!���L����<�=|q�i�,���v��G��"���P^�P�`�s ���6��!���7� b�j4�dE+����B�� y�(G�;e>����!��6�c��i{��W�FW3�#b�I㬆�6%zL\��*X�߆{ۘZD��#Ry��m���9��.���瀠�E6�q�#�(��U.y8�����b
���e�o�_��ek�)9�����@M2W.-��-�4���������i�L?˅�����~ڸ]I"�"��^�Jh�֛�����$����Kçh�dw2 �i��宱x���.7�n�-B��45��5��BI;%S�@%d������R��t�I�����̘�iF��4y|�02��qn;�\ǅ���e)���
��d)�����@�ً}�)((�����W��.3�6�Ƶ��T��f��X�t��c�N���k?�NE�C`��٧G�3��<ެ��ūd!�2�Ms��[,�q�!�"��^t%$��K��=�u�y"�k���1(˧�����c1[w{�|�0	�}��o��!�9#\.׵�ږV�@-�'����~o	8���yp��"fZ��j0d�O�[�9�c���O��&U|czPǥ���$}��Dֵ�8�t��5�FM�{]�|����nT�sp�o�r�(��N/��h��>���2������w���c�.@Q�֭,�`y'��TW�ʱ�2NL���B�������N��!2�!��0u8�ȥ��*%���)��h��y"�"�F�[�QM{���Q#O ��2 ܁����xY���t�O/+���8�b�-7��\Y�)d;���f�YQ*��<��(^6Q=�I�������93$�IWs�}1w&�a���w�㤤�����yY��}���W���ʼ����T��|R���t(ה�
������AgEh�]{��G�A����d}b��d'������w���̿��ݟVf�ʮ���k3Ŏ	H��Q�w�\H�x�)�u0`���%y��Ek���=ˬ~����+�b���4(>M馭�׵Ȇ��� T��'����� �;�Y�*�:�oh�h��������du���Nqv3��L��Gk�J��"��3�b�|'|�~�[�q�����l(�]9 \mc7%�����������҇��~#גbC5�O�!��o�PT,j�T�f���\��'ß��E����מ��ޏI�Rɾ9t��,�R�5��@7� �\T��65S�C���ٚ��C���ee�6j���Xhd}dQ&A��^���n�I�W��QM%�w#���A��|�W������:�D�g�O�3�Z-�y�8d-L���2:a�w�$��[�oU���V�nfϘC'{'�oA1k#���]���|��چ��&p�.��^AZ�m�Jz�{��_Gܮ�O��GE�j�.P�hf_R��.�ք-�1ơNOD�X�/����K4�@hd��胨��ס��T?+��Y�B��;��O�-����i��+A�ɞ��(�P��{��	��%s�c{��7���ay`�U�WiG;��9��%~�"n�B��")�����V�ǝ;DWttހv�]���u[DIm,��U8�qc���i����-�ׅˋ��-�@�W���\�ȿ��vv�Z|Я'<���si�-�#aS��Q��v���UF��2���7m(qj�q�Pe�iwp
�𜮠5���RqJ;@�����,�"&����&g V��g�gg�>P/`��t�bt�Ѕ:80�fǕ�`����i�r�E��W��(��,�S�h2�v

���n�����G��d�hW�Å�xb�=�/e�:v=`0\�xǟ}�3=8^o\�ʉ��e�aB���=ʔ�5����͆��,�*��M�=�l!�=S�l*0fLpY��|~M�^tL&�/ܷ�QP�d�DT��<D�Ũ��b�T���⢭���0���)��\�I��R�{_�}�7�q����Y�/G>����D�2G��2��RBt�m D]���Sz��NZ��97�,�,���;�;�[*yR�Z/��.="7 |�B�ƶ�T�v���Ν�gW��*ZA���=C{�G�r����s��޼�8b䔡	�X�K��4P�_��.����R��M�?����m�~�F��:eL�b����Gj�8d*܉T���su��2t��Hu|�G�umr��ؗ��A�;���?u������|Ppgr��H�+��
��r߄}��3���8]��}yDU �p)ƒ&ٓ��n���X����� ��k�e/v��5�x3HC��9��e�J�-�<�����~7:��x�R�����RU^AlL�v[�;���F}Q�����!��JnՌ��^�.W�I�f���_.�5=�K�=Þ,t�{�U��t�)��,�� r#�O���Z�U0mB�8;<G� ��]گ���{�Z6�Ś7q�,�k�܉\���c��Ű2gDf��c��t���j�4�D������"����*�E�D+��d������+�"(��	t�,݉����a1!��-+G0�z�|�
�r�A�S�i��@g��?�-����Ӥ����m��[����c�����W?*�d2���M���u���x��݋E�E���U�{3���E��R�G�8q��@�JEQ��!�X=��/�ct�b�����d�G%�^ڼ2n��T"�B��rDG	r��Cb���xx��F���khZ��	 ���
��Kg*<s���'�Í�m���x��$���������na�Ȝ��'���T� Upf(��%sعnuke����;�x��g2u��#V5���,Û�yay �EV���X�1"�	(w(�{[�Ԟe�X�
���s1P'�_Gů�7x���T��я���S8�V�� m�:��nف,�R^��!�d,V�,�ƚ�!���ic���e�܏˘Ð1�ښ�b5R�Ir������x�,9J�1wZ�9l);���Ճ�jyo,��ƘQ!L���m7>���e�j�s��_i�{�ͪ���Ai��d5�\�*���Hp�����l*;$�"t��t�I���`��/�hס���i�=1Ŋ����m��kkio���/�y>@�}����⒢ &�.��W=���Z�����2��SNM��(�#�^���]F]N��LU��»D%��ɇn<�b=u��c�^�DsU�>&�f)��w?36b�`mԄq�I�����}��e7� ��4"�BMA}.ŝ��p5-�Dc�����c	�t�\�Q�)mN8�/7���5�r�p[7V8��][u�e��8p��ڃsϸ
��t�K֎��T�/��^�x�z/��"
��]�t������*naڮ�s��Mj��B���8����n���tv��Z��P8�	sT��<���Ikځ�o_�D�9#TQ$�����c�Ö��255A� `���V��BL��ː�rM�R�S���F�J&�E�,��/�� �>�N�l��kT�!����e����&jN@܋f�/$bED ��[,Ӽz^|��4��Uw#|m�5��Z���Z�/��x&Б?�,}$�J^��^I.�H���]�AM�o�F�Q�u�:p|����v!vh��4��hZ�5ı*� ���'�ȶ1�cRJ9iErʼ�)����O�)��
���m��Se�$\|R�uZ��ñ!�Ǔ����ς�W�_4D����ׯSпﻁp�%+ߣ^Yt�����U혧.�sh�
����tg� ��a<^>00Y��!��<�Wy��2���v�U�ڨJ'^��p���[08�����������e<�}�:u���"i�	.��c�$|����`؉���EA�B����[�h	�a�H��Y����̰��.���p�K�M�|r�W�q�K��*~����Z�śbڡ��+�tB5�T Z9�Zz���ұ��/�*h���`�K3���]���������m�����a��qA�������J�
��T;56|�%�k���j��7��F"�ޭy�Q����.|ǉ�홱
��͗�A���]�$�A Z�(�c-9\��W����v����A�a���؉��LY̴�C��C���<0pmK`{�{�[���������Gg#�3�A�d�s�}(��&�=S4Xb���/Q-Q��̬oZ�p<R7C(�V���~���p���L��:�>w���l۰�;N@� 8n��Z��{Ө��<'qE�����+L\��q��-���A_|�F�hИ��9�U���Et������|���1�It��#F�[�c�u�f��u�dDޭ8-jD�	��"[��U�mf��� �.nX�Fa�foIA"�LOCr�V�	V�J�����{������ӆ���o��*�o��vC�:��/z��fg,��q�fP�s�r}iy[0�Ft5>��iS�WY��L�h]�?W��գ�_Αh.<DB��]�yX_O�Z�}Y�7��[U����j�5�gv����]ݻgJP��84�����D�WCzb����73ۼYQ��T>�=
po\��_h0.Xz5l�f(ek`���Zs:1�L�xI��ot�5�t���YO>���[�K	dꎪUO�j�զ����f��IQ�q;k�䠆c�-�y�8���䁪��Q�7Ow���T����E�8[���A	?;j����!�+��1�� �R���1nt11�Ex8h��x`n����=U�����o���,�uڏ��BRR�94�tSk�r��� �<�ql��ې�q�[N$��������}��XOtB�T4c�1�8��C��G��8�1���+m�[������o=%�L�_��ߦ?�6��M����&nԍ���G�+_�����v�M���]�=i �s��:k�=��uq���gP��9��,�${�Æc�lQcs���
�}/�yt�'�x���Pk�@���R��TQʳ��N��֏c�b���3W���)x����E����%ZV�Z�C_��Tw��5���sj¹�ql���[�tB��X���vf��(�A'�(.�C�2�RL}�\6�����Y��A�E�0�c٣@jS���4��k���6�������x�P�F�Nु��QB�a���cFx��7|{��[��*�O�?��G4ɶ2�b3�C5�EI�=#{:�*~p��~�p�-`����ZԽ�t��|�	K��p����ԛHg�|A����v�$�&q�y�4pH��������4Nx0D�?��!��(tX݈��^��p~`i�iaix���U��~
"V�d�S@ۻ����>��񥗁��2�wr���'� u����VV�߆-n��Q�X�̫�
ܱ�n8�tФ/�o���j�P��THJ�� ~�YD��vU�J~�\�O��ֶc������=��0ت2z��Q&��e<�׏�,��P��JVSC��[㻅�_&Z�i�E�{o�|&-̆�_恁�
Ɵ8p��#�N
�h2�C�n�K�͓Z�7���!�8��@]"�Af,+�%?7��A\��aA�l��VBJ�����q��w��F`��V�0��x���^n�b�E�M��ofw5�ۏ���䯬i��5Ҩo����Qc�%#7��we���������i]!h[�ޮD|'����ە�R倉�.8�b��O��1�̇��&Q��);�$h?��ܲd!�DV�p���Mf�d�~٧�ϑĉ�2;���,dOj�����Z�����r���MYRN�]P��d�ϵ��xm�Ҙ�2��U ��^����{]��o�	i��]���kj��d¾�2i��VW{7e�&�iȱHDT�lg�-��ꎖ��bGA���w$J0q��,?�:p�������*&D��/"�d៺��"L�� ��c6K$!(�D5�|����c^�n����V� �R������:bko�u�@�N��/^�r�4��g'�:��v�/�%���0��{s&P	(*����#�#>۱�'g���|#���Ȧ����v�D��A<�H)�`G�C`UfcUaӝ�kG�4�te��� SDūR;�� +����2�"��&�����eXW�d�!x[�7�`E��n���`*�%��=��-�p�R�uWJ8�G���{2)�m�5���9�+�FIz��Y5���9^��rc��d7��������|�D8Q��+q�5T:�7����T΍]oSlh�h�A*���,a����Z�����2���\� K��m��E����e֥�Uߋ����1��~1�ж��i����A�5�[������W��kI��V4̃E�X6��?���[g�"��
"�7���\�7xd���<T��b��R�\+����O�v�'���l��E;x�)�y��c�kB�/����bG���_���{aўN�����gd
�f",|��z�9R��˃Fz_B����Q���4� �? ���O�ϓ����o�JՐ��mK�e����:_~�Z�!U�Bz�BsT���#4r�H����َ�39rz����O��a�G�����}Y��=cQ��nAp�?aD^E�Fq��]�
g��x����Ry C�>1e�BWT��2�1��T����`�(mJEr.�JC�]8���N���4 ��j����<��Ⱦߺ�a)��p�t'wnE��9�><��e]lQι��F����lau�zZ�n�)�PQ�nT�����i�5����ź�ު�$JY!U���SX����pu���Tyr��{'=��y�7i#/9���(�ES��;l�j���FÙ��o��I%ں��Kg5�2k�JI�ZS�(��d�y5� �,��T11�-l�Ϫ��=q|T>$Jw�O�ihӵ��.�3�Fm�`�Į��ߢS���	=[|t�b	VɷW+#9��㠫�W����!;�	�p�y���d�9�.�z�'}MՈ��Ws���$���[��)�5� �cvȜ�K�#��vvic`�Lm�.��O�l�'�z^�NZ������6���� ��Z�-!���~���^�ɫ8�zL(͟�V��Z��J=�)�����ۤ��M�rdzGWz�������{���f^��7���7���J ��fGq��?)M���]���!��Y�̶�%�ہym��y��A�͜��c��P5��	f������5|�!^\T���v,�OTҠ�w�q��o�0�����xX���wETe!_��@�A��J��C��d[�"����6���Yt�he���m���^�	���,��B\sI�1L�P��=�H���}q	T'��l�Ie�k��>/?�2?��qQ� x��3W��Z*I^MZa뜙0	�ş-��ߡ ���^u�)h}0� ���R�"�Re���%LƒB���a�^�E1�.����V�G5����CiU�pQϤ�������]3X���y�%3�|��Q8�sU��\�
&��`�����=��z�L6���bl�s���wPG�Δ������1I�qt�J�(�7��hW�\�nM[g��fF͕����(o��0�(-�ڠ�r=2�Q,�I(�Y𗀧{��o�

e�#�a�����'���i��*��YV���{��i`�C���ܟj���Z�4�#�~�d~f�
e��;��p�p�� vC̚�F�t:@.$�������J�^�	uC��С��cƺ)^)AR�>����
K�_���^����/h�����+N�`r�^���I9�'��~6��M������c
�6E�NҠJc�}�a_���<�i�H!�4����>�M��h�y>A�c�r_'aw��2��#D���k}�J!+Y��>��D��X�(z=1u�knQ�1;�4�p����3롲,J��k��ۙ/\˸q+Z4i=3%�*KQ�m����7p�%�#��n��fCl����
�d|�nD>@���v��5��	[���B1�Fh�a^F����%E�)��1C�{���1��j�>bAʕ��|Π2<����rF�h\��e�J -�'3�_=��&���M�>��b+dc��1b7w��r[�wm-yj���O��C��W@�~z�|F9 �gH��k���ȡ=O����G7�YwJ�X���Y�}Ԛ,���9����-,��秋�P��� $l����#��+��a�>^�~,ҕ(�Hf�~D��Yi�T+�ߍ|�~�	k��µ�~�'nR��ɥ�JEi�}��	߆��y��{���B��Q�)�f�wH�a����Y���t���/T�On��f��Q!��CK��Wt)�i�Yt�FwU�ʉ��Z��iag7���xMQ�����Z�RU��2h�|x��F@3�~<���Ұ�Q�6��,dܶ�b�����ߍ�=�m��N�F�ƕ���':Uh+��G�}�g�9/�q�DK;9G.�p�o�zj���8M-5]��/�&y���Pe��_լG:y�8}���(�h�8��^#h�{a[rSd�j�I�΃�m*,��������`v���@��� 6B��DDx��j��p�\���6��{�S��0f��k	p��|�Fm�=/L�!��9�ias��na����wo�7����s�u�Y�������u��n�e�Y.y+[5-m4�$�MF�v��l���~]=�Q��ˁ^�" q�����|���D��,zhq�&��������-���r��#g�seHhF5�ƍ'�V��#%P���-��ƞ�� �}3!�)��Y�D�6��ұH/�V��>HGh$B�P�?S�B.-<��&��C����&���}Gk�1�?F,�b��LxĠ��b.� ��t;��Z��L9x��{_c��ޝa��YJ0k���>kDxd�i�٭u�KeU
�%�q��YA���p:M��\@�O�v8���'FC�ӭJ�9O~�����Z�A����q&6��-�נ��@t /��т�p�A�>v�^{}�d[�cwmN����{�Rn>�0��w�n��F���Ě�����E̋R�/?�f����CiZ�|\�7��ClN�`w(O'�3c�_��bU�˫�s��Ɖ�l/�2Ql'Y<n(�1���~F@����q �Ku���Е�J��&�Ɍ!Se&[iS?�60���i�jcc�<�7y݃�EY��ݾ�j�@��)�9���J������A�g�/$���5_b{MKR7y9_W���Q��vJm�_���?�/P��5"o�dK��������D�YeQ1�J-��?�73����Q��!*A��A$1- ��h6;u�����t��Bt�Vn�����#�<��(j ��/�<x�Z��lz���i��� gGG9��B�>q��\�#o�1�~19	i]:��B�?�?��"8R����GK41>>�"���dx�E�^�v�@�i?l�;�`+�8#��ɜ"��0��X�8P��Ơ^����A�Aĉ=3� �$���IР= N�	$TTm.�����6���<�c�L�����ɖ���V�TE�F'75E��Q��{t�߱|�|�K������ϼ�0����� AQ�%�!���\)�dF}S*R������t��DY/����}%��!���k��|�|��ͤ�]��R���f݋�I@��-5l���Sb$�;S*O�G�����k�����|����4J�I4|a��"TyALy���
1�($+�Y��@'��#�'�@6Î�L��ᵃ��&����U:܍����̌P��
�>��jp2#K}��$�o�|hK}�/#�v�7t�� %��I67�����2 �p��I^1ھ�Ke���[Fb9�ܹ��ic;z"�d���?C����Cz�&D�Z���Q�Y�\B�:�+SO
��p�_��o�3�n�V3��)�of�	���`@ZMٟ�O}���ô�&K�oX�z�p��F������XѵFC��JE�䤪U�R�&T��to���
�=Ȱ��цM|;�Ǉ{9��i~~�>�H}�{&�Kw�!K���Pk�%濬~?� +��J\C>�������fq1�N}3K���x�{m׻�Z�G)hlZ�(�7̽~�-�ø�!�gh�2�c+B^*�^����JLd��n�*�Z���H�,��<�p�N$����o�┺�%�O��tʸ��0E�%��}�߼}X�Z[��}��-���e3��	6��� B���"k��+��^*�l������g��0�����/���)�w�.� ����vq��d2o���_��1�Ćj8).u���6A��qWZ���k Ϭ�ͪ�y�]�w���)�t�/R�N+=.�3[Ʉ�h�X;��z9!��������>r��h$J�� 0Gs�bO.�:{�?�º�52�h�MW{54��mZVF��'��î�-'�f�T�M��x��6򛢎$�[Ua�� U�dbx�v�
�,>:ꂟ���A4>B�q`����K����z���3�Q��3�!p7`��K��.u�\RRJ=�
�I8~+�3�� ����3��^`���M���F6(�w�R��E�t�C�<�}�N<�2d�q�.nȶр�[�Q�%�& ���N!m�I��/|�R'�������"��N����^LC��^ŷb�C�Q��GΕ^z0��2ϯ�I
�م3!m�	�
1�C��/�Ә��ڢ���� 	>��Չ����[��B4#�Cf�|���V�����R�jɶN�D�?[[Hq���+oBBA�gCHPK�+^����CU��,���x���c%֮��9��V� )蕶3���̜9��M���$�v\�0<}�A�K��Q��A�v�� -��u��z�Z�c[�pu��N�'c$\�*	���HA��������K��f�e^���ԟS����-<<�3s�����9��R<����:3-��y���f��^&���Ҥ�3�|�,�f�<G"����.�E7D2@�|���kU����#!��(0�9�ܶ��4q�XY�e�ת+�ņ��������+*��Y��eP���ZZpѾ�;-�Q:��|�����А&Ԟ7�#��5ѯ&ˈ�[-�t��'��Y��f9߽Gw@gR�򛖻��$}��/	I��<P+m8g�6P�A!,O�5L�3��|�f�����)ΐVײ���s�� \�S���顏.��w�z9%���>�mbǇTb��Ur��dIۃ�?�,p��������;<�֩��X<�ٯV'(�!	wh#�����p /K��1(D�-V9�Q��vuRĕ��I_g�K����v�db�`Ӱ�3�F�)my� ��0������Fo�:~�}J�T����g�K�yB���FfF�0 ��{�vz�J��	~(�P!M��?��~}ۥDY:�7(��l��ۻ�Q���� 4n,M=	b�Bd 19e�M��T���na\�٦64�<�~F������a����|Q)��MYZ����a�+S���r,N�c�r)҉I�\��dg�L��<Ѓ�	k�����4��(s"���]�z��DPZ�hzS���u�?G
A���QM[�O���`jۊ������w�@���'K8���}Li���3��t$� ˕fA?�}E����T�$4���Cy��Rl�D���6�fa^:i1�d�����=���k~n�%��p���8�E�I��h둮�O��8��.�F���<Elx�� ������d�a�S���I,��ou8m��� �Gؼ�c���'$��[-$�rm|A�ҭ{�B��=*v��ث��p�ax�w��`�Q�/�xh٨H�ݗ�J�Q�H�C�B1V�Oݰܬ/,p�u����q�Ӑ@����K����D�Q�������c��r�H��S՗�H�:����ҏ�@�^(i���2��P�} ���E��.�j�T���l�Z���;��s�\�����AHa����3�7K�� ,wK��c�RW^1��o�ώi<w��{�$�OJ�KBH�7����C��eh�2�ΐ,�����<i�x�Lۖ%�7��.'j��F㘣���di��Ơ��Ka����h��vt�?:凥QT��S�}l�_/�Y����Q�M�N�N�]F���T4�+E�HiJ;���D�5g E3�j(K����@�w��}���i�l՚Sp.�C����h��X�>�_�{S) �a:�	m��G��8�b�a��o��?�E*=��i�ʀ����\xK�hF*�5"�@N���[N������	���=�$n�+�ś>�W���PPVx��_Y�o���"�G>�LzN��mYݕW��,�3j��9�:9��Pm�/���
������c����Y2�U�g
�B ɐR!S�A3�'iU�2v ���J�N�9")��[�W�[}m�_\�`+�6�$]~`�"ʇH��k���<+�4�+r���(~��P�,P�=���l��}'�\DYi���(�_č�m1]�D�y�y�B|v���|$
ě����pU-�O�@��L��-2_o��ۆ9�_D�}X(^�zn� � Lx&�e��:��Rn�Z�g�B�u��u��XZ�������;w!�r�9~��n���6�r�{�:����P<G]�	��!��� �����a�L�.9�E���L-O��� X}��U�-��(:�F�����ep0�x����{��8�|��:��$�<���88��N�Lr���"i5[��>s,�������ϳ&^�i�O�B��Ԅ�-XF+���~]�=0�5���#k�g5��"�Jl��䈞0{ťK$�q������r7
e�Z7"d��X���ø\��j���� #*���t�ݰ ��l8��$\2L;@��v���In��M�h)�+�C�^ď��''�!P�dtx�Oހ��>��Q���O<���6���@%
��JM �)��܆��q��t ��N��j~Mʉ��F}�=\0��T�}ζW������F��A{;~B^��H&�L�˲�k��:�>L���8N;�9�.���~�,��x�������`tBU׈�*#�v�.�ڋ�˳��ҫ{#�E_�E����̀�'��n7;ҕ�iˇPǝ�8fǂk�N�RG,/�b��˂���|��I�8s��0s[â�V3u���T=W�W:��֫�e)�u�n'�ׁ[�![
�"rk�����ZId�v�-���&#ٵ���P�ӝ�Ե IR�o&����t<�M_���D�Ӵ��q���K�n�\2,�D�
{a}�3����[�Y[�Sa���*�@#O	����V!/�C�\U��;��5%���}��� 4����;Q �]j���� Ħ��`� V�����r2�&��2g;,@ǣW�z$Pm'�=�����z����>ɶ�A,��~2	7N[�5O�t*���-A�瑾��:��������1쿲SE��Sֈ����+��av��W\�<_��R�g4�ˎX�w<P9��Ġ���j"�	ޤ���7q��u��6L��ɟG9�H����F�{��[���&�<[�eNXF�Ce��ζ{�D�Q���c��,���P�P�Gqf/�x���IrWW,��_��=	ߏ��}/�¨V��!���<�2��bhYK
'�M��{R "=@�cw��ބ]��Җ����M�'�nǾ<��Ӝ���R1~ԺI�=��CQ4����E�-rO�k�X�&̇��9/q�/d(�lN �_zR@L�'#�njy5O�����P�YS����7"t�S~C̵yM���D��;i�/{b�{1�L���w|F�."5Gl��w���r�� ���<_���J�c�G�o����*�r��X��<޵�����U�~���0x�ګ0�<�K��Zw�TJ���|K攷`)�����
`��)P�qϑF�]�!u%�D�Č'��'|�C�+M�����n6ϛ�$В��혻�v<��+�������H"dP���A�s=� `}&���G�.A�������HP��T�7�ẅ���E�6�K1=��}������ٷ�)<�GzR��b��,�C�M�)��n�`�<�0)�E���7XsK�m�O��ԒB4!1�}���Oq��QO��!��Й�3K8?M�	W���B+<���ծ<�ɞDQE�
�s�K�2�u��j���p%�W�����ڹ�*���OR��"�%	��B�G�,�A�#e��Y�� -�O�(�Q��6�x�h�5d�m#�oz%L?��_	Z���ug ��D�A�c�)���� !���~:յ���iuJ�{��K���a�0�n�E�*�#	�5q��w*C���iԂ�������`�%՝}��՞�'�
��#J���,;j'���>D���/�>ԣ��Hu^Q��ڝ��`��E0�y/l �5��)����b���tcx�B��S�iU�Q^K.`�-4�=m`�0	�����*l�lC�w6�����[��\@�`ܾ+sK���W�ٖ'�!�n 5�PT�����յ�=U�.e��	{D�}3��Nl������&UU4�%��a�w����	((��e���:�C�ӆ�.��2gqu��k��i>jn������T,(L���h&���8��{	Ʌ��ިꌊ�+�����o@k�<.��	+|�{�B<=���<λ*�"V���F5�s�mSn����rA�x6 ]9��	}Q3.)s�v�j���s��X�J����7�XL!ƞ3���K�X6j��OƐJbO� h�"
2��x2�'��,��9�9�M�U)���*��j�g�	��M��Tmv�l8�W�B��[?"b��`�)��9��΍#�\6��(u	�N��7E��[ʠ�o�!n��
h�3"�3t�������Ψ+�Ԟt�'�0<��A8�ja|�C��]�7v����j��I4
������ 5	� �i����ם���E�����W�F�ַ�1�½24So�������F�d�	�y�,E��hK��L0��܃1����si�o��pոP79J�7��U�,�<r�<**	*�
�pifm	�^�c���r^0�?ls0��u]Q�y|����
"(!�Z�*�G��(�E��J����b��#���ŁA{�� �"k�I-s��pHz�l� AΝA2�,DK�^r=Z�~�q��
`�jT������"�H@K�'��m�C�
6��~�c2)�sL�\ԙ?������?���P�D�n��W��Ⴝ��ߏ*�Dc��l<���e*H��{���W��B��Ra����P�jۯ����[�-�LP���W2�V�;f.�Je��f"�kY��%����9�@ ב�؟���)S���0�?��*�Yf��҇�g-	��� �=ᘤS)؀K���.ec��j�6���[�y]��k��'K$�H}WU*��ΣEn����\u��M"���j}�O�x|�>�l�I6ﹱ<�L�Bm�(���G��k��~�.��VF,!#�T��>E2���cI_��|e[�AR]9�R_ؽdEQ]��C�2A���}sb��Av�m&s ���G �
���H�=zi��=�o���]
�t8fj|0rPt�Hl�;��p�w>�ۜow�|�-9h�
Y�8x���u�)��(�P=d�:߄�B������<};�U��>��jS�e�^GE��d�m�ˍx�Z�4iY׀�T���6���}���Z�Ͽ�Fzj��%�esdEi�\��ul�5��V��6�]=�N�M���_�
)��QE�G�P�i0��>^zk��f��_C�N����_�-L�8R���o�`S�f��-q�8�ZK��o�<41�U���&H �;�m�qˎ�.�fL�����W|�f�~S8�4O~�00�}R��bR���4n��OL`�e�a�D<��|w1=ۚ������&�8����R��E�l�'��fSSh����g>Dڇ�rC�nLwFƿ�E�LH�Wf���ge��y�G�ny-�0{M<�)���J��k�L'��6z��`4�c*J;����r�M*�+:�����N�n�!��4$"�֍#9���ĶKO6��q9�N2��@�B��,���5��{x�=���bO$�k!��X�|8��H��.�8;�l'�C���q�B��,�l+\!W���\���.	�
��8�пW�E>��uC'�٘�ڞ-��Z��W[X��o�L�y��]4��eyB|���D��3 b��:����n:�;fgk0����~
s�
�]t	��O��x�~&�U[l\�=�m�2�������~Ԝ�AP4$y,�{*�o�	�kR�U�k-d���&�����N�v[H2w9ք�lx0���d����2q�1剕�ճ�v򮡾�""��̼����e_�eK���c�Ǘ�]� ��X����Pr�vdǰe��B4�^�/d�O?�1;s�@��X0�t�&e��"�-8����0���(�B6�i<E1��E�'����*a`b`����8+�7��'=:�*�3�� ���@���-ܳ=FH��0M���n<̺��[��֙��ln��1m�2���(#4V�ǍvB@Leط�\��/�#t��g��t7�#����BNm{ N��x)�4�
�73�:p=&l;Cj|�yG.FKi�nJC1���X�D]#haha1ݐ6z�Ͻ�>�g��i�i^��CpFg/�'NR3�F�#rPBW��J)��G!L�:^YT���}G����*34sUw�����\���м���C]W9=��eش���N�8^X�K���2mnzM�����V��wR���'�"����k�7�P*2����-O�͔[Q��9k{y��X�x�A�~1K�����A�N|!��Y�~�mkyn�lRyH��dt5�;��D#�ЫzAjť+������s�:�[�W���ץ�i�u��o]2 ��8�ͩ �8�1���Ѽ,s74�i"5��TX���d
R��U�-R��(�V��U|�3$Y\�3��C���e�#��Q�}X�i���k{��_�I/g�<a���L���98	��t!���6IQ�u�SV�T�f�U��͠W�����I���Щr������G,��B�=ݏ>ٟ-S�$��TaX,A�'b�,��^낐�C���A�b�����X*������N{K�lSp���c�2�)���j�o|F)*%��D0��y{V�s��(��w��^�:O��^Ծj�&ba�S����������DBc9��c�7���
&t.l�٬�j���[����Z:��?��G;�iԑ눨�aNJ������9�~K�Y5�N�,	��u2��%���.�@k����]���/筂/؁[nd���X�/����y;��;�ꮳ�.G>�2�q#i��L���,��j��s[����Q��X���>�\���|���@�	Y��G�G7N���86rs�;KF�LB������n�9��^X����.yc8�2�
���	���V���i��H���Ҍ�4���%`e{%�buI�ٽ{�	%�A��p���p~�.���bbi ��b2��S�2�̓��7S8Ъ<�^kɆ�Ϲ���Y�����A�x�C�W�t�J��g�v-K�S�V3'�0B-w�u}�@�.�XZ��9`4�?y�<��c�
�ۭ��<'5~<���~!�aڙ�r
�}�� !���j�$2���sRvS(8$j9��]s5���L ��w��d�N1K��X~��U�H42�� õ	���~��m�*iր��9���JM���e�'g�\ȱ9&�K�`{(,XFr_zI1�	��5U�/��Am~I'~S�H����6��?`)�m�t�Ė�2>�r�K&V�"O�'�I�V�@��]/�s� ���q ��b��c����~�k���G���ضv�w>��^L��u&�(�YP�
�ȡK��t�7��-��t�t��&d��N��,N.��*��E��,��ש��j�3��:�`Y~�d�-���;ľ�ت���Cs:/��q|t����l���"}Óc�f�Kɱ`n6�o�#�j$�O���/���>L��,I���b/[I�ۀ�m��>��F��C��r)  �����،��߳�U�O�ihQ���i��E�*Lr��6�q�T�+ ��R@]{�m$G��0iܭ��Ԃ.�=�_|�J7S(_f�H&j�f^/Z�,a(�cOV�S\��Ο_\����f��鈟���1K�;�z�eٌQ�,not���wb�����y��|�0���	��U6i��%��To+�������K谝�ú�����%�ZG�g�e_����e���cn#T���娾C1���a�Gҋ^u�/:�֨���W�y�OMJ����Hlt��0�#��1&Y3V����I�(X���B�<�R,Uw���U?��d��3x<r��8�f�˝��J\~�:�)�()(�bW��*=>���l�^�NξwIl�d����}Y:�Ә�L'�.&��*�� [s�C�� [b+�_ _�.�Ұ�5ܱ�۪|����ɲ�KC�
�IA���⥨s��99(���|�o�jm�?~YW��d����C�c�+�����$�V#x28X�W�[��ē<�3:s�۟��g�q�>s?Pp�M4�vh�Q���6��H��+�	�fȿ���K��� �Q�܄76��N�Л�*��}$Y�K|�ctA'�����$^��ZO;�4č��Ѻ�GO�֋v�7�.�?��.��0��]�Ws⋮��+GøCf:M�W��"y�vY-���Z��!��ba�����򹔴ޖS��r�X�J�fj`-�X�DˏB.��`}��-��,�EnD��Q�{��S�u��������E�@˾�	ȟ�2�)2ɜ�}:�� �t���DЧ�s�7yim�fE�$Q1���h��!8�PƁ�����%'�}����k����'��^f�]��!�Z�{��S
U����UϚ�<nl|��Y���:���x��;i�y0%�J�[4���/��*��K�?�����깦3�&�_r쀕 ���I����>���+�����%r�  ��f����/&��!5�W����@䑠!@��G�IoN�b`@��X����D�:����M�n�I)����e�����`h�F�!+G���`+��E���*]}6��$��2�A�K� ��ᜋ������͌�Ʈ�2�=�':1v���-����{|���J�B)-˩�ԥ1(�@@�b��R^a�v+D&8����gȆ�����R�W�:W�]T��/��F\�,��R��''or$��K��W���fz��e�nj���C�.c$ENi	^[��4�#��Y��V����Y`1�C�3�Pp�%�&��(2��� F�m���e21�L;�@$$��a�5�P?�rW��m�p h�u䊙�����ѿJ͜Mm|��Y!7��K8L �}�a�2T%x��(�D��k��f&�O��P��(-�F�k���/����nCS��@[.�_&Ju�)���YsmĒ���K��c����������c ���h����q�z��|�t��J��.��۾�t����y��)�p+�|�̺�a@n+�yG�M<����ϸoy�q���x08]�v/m�ti���JMk�)Ŧ�)�J���umV\������Co+���޸�K����I��<r����ZtI��J@��� �[����oq����o�F{�F�������Q���Ach�:ʿt@�֭x����# ~�wI����עK��
����4�i%�h-I�������ɳu�͕b��p����(�s^���K�� /P��]
�/�X��o����}#M�,�eBzv[ɹ ����C�/D�\I_���kh`��&�Dt���l�D˝]�Hr���:��	����ꬮ\g��'G�BcY�(U���6�ݗ'�~�7�F?��d����C:a������z�d*yo*��*W��΄3�t!�~_	*5�~֪����&x�o�h0�r�w�D����/	\Ⱨ0�cs�)*��7͉xN�_���V�}�{�������j��7�I�)�3x������Qngb2�1�p�\r�\ĮS���W�G��s&�$�����/<�uF-�ġB	nr�&Щ��e/v�G�����!Q��}�#�;���;�7�*6�����Jo-� �c3f���Ms�`�ޗK��_�O�aD�*�k^�]氾��9�"�{��4㚆��0ֆ�ME;�<O?\#��l�ҘM��ث�����J���Ǌ?TA�@�ଷ�D\� �ID����hSv��?�g叠�I�ms��qWz;i�oR6c��7�My����k ^������z^S�-���6{E���o�����(�����SK��Y��v��!X�s�x߱����!�Ϡ�F�XVW��CD΂�̧m�$����MuUc%�f�-릋Y&얟�$�-��f��w��<�qiB���������-��sg#���P�tJ�r�����>������ �������)��
&]ܦ�:��#4O�o�­���b#��B�"r�JeRBr�r0 ���Á;�7Ijm�s>g�f-F�
��댤�\d 9�:�s���T���������/�Z��m��w@3���0ܮ{�ň��zt��3'���`�����Q�j�� �PJ"��T������o1*k����h��#�М����	�z�R�.�A�1�a�J)���s��V	?�h݋��y ��=�F��{��ȥ��Ej�o�)%N���/PƜ��KA��ďI���p��+z��?�`�8��m��ɧ�c2$���p3�o��m�67jG^-���	�m:������)BO/.����Z|2�N���9#��	� ٪���G1�\��2WΪ̂Fc�OA�R�U	~|-��f1�=��T&�b�w���舧7��3�������J�v��t�6?�z9y��x�miv�����UQ��4�/s��ID&�W:��Q�QnX�$s�˩��pί�)��W��p̬�A*�-���"Wx�����t)d�g�?�U��b����7���/.��?4����]�6J+���4���Ό/�p	$3ۮ�.(~"��4����+h�(W�3���ߜ�;��s:���7|�Q����;���c\��s��	��L�G@y���p��eA�L�g�HA�2�o��f���/}LQ�/7,p��v�j�S�5~�}I4�l�q3m�y��!������)C���Do��#�J�.�g����Y�7�����ի^��Yv[��0{ؤ~^�,%�?��T!��'��rH���BJY�<W�7�����'tv�8z�����l�G:���J�{���V�`����QY炩Ұ�-:�;G�i%>�1P�5"���P5�ؓ�>��ax[�?0n���_��~�������T����6���:���=���~3��M��!ot�"_v��� [�+�{A�ߴj8Ta �PX�[H�l��xJMI�c�b��Ew��5���K�/#K�Ύxy�f��I��gσ
���!4̐&���MX?Մ
��S�k������њ�D�Ft|���4�אP���K����8�˙������6�Nx�4[�sҞ4�"�a��"9��B�Q2V���-u?u�^d��ؓjN��,A1���#�4��M��;��vHJ�5�}��a�2��3�h�h��jR���Ԇ�4q���M^4�����H�be�?o��U��d9p����?B�8F>����/�zq�6�C�<{�,����z��W�tB_���z`�����Yiz�|^/ �#�)IZ�^v9�jQ<Ńd������z-����Ը��S�K�&�"�� d����T���oD6y�O�����{ة <'.��+W���	pDH	XFs��p	���7�Qyc�U
��H�}���͔/ġ:��G�ph�BBQ5��	��w�=����)^�xS�&A5׎�K#��}�'�H@;;��f9N,��z$�h��K�e�Y�K>%�O�$�Yi�L< �9�����]�u<\t ���ʹ㩳�v�~`r���`��-�I�m㺥Ϭ�!Z��󘌠U.M���陆[@��/�Rݘ�;|��<a<��1��{T�N�֒w��˄m���2�@��{���jd}�q�&����t�������u:�*/����kԖG���^�
6U��%����Ӗ�u�@�ɐ�`?����$��y���)���+��e,M�yM�x���M$�aJ���kh"E�$��E����F!S�/���H&�wS;���6$�_��_<Zn��0�q�0%�=��� %��U:���9e)�91l���WS���SHJ%��s/ˊ�~����=~���|�,�nK3k�(c���)�����&��tt��Z'LX?�^�Q O4u�J����c�����0�	jS>����To�4v��ɇ��+�IȰ�O}5�3�x�*��-�f��I���Ʃ�{Lpl��<�!H�K"���̈́�1Eꊋ$�>>�o�|�hV�O,��H�۷TN�����#���8/g���J3���W� �\ݢ�!�_� q�
��MG�?=h���O4~w�56�3���A��:n�%A�R�?VuK��L܍>n�#��h�,�p-���Lq�+�U���Đ3&�\�X��
 {榵���;м�P�����J�4a�M\�h���*�?g? w]~�*���+Ds�E�=4?�E�%^�T��#�JrH�
,3`�_) �_8�&�A˛�Q�6�����+n-<�
B~�EzbNJ�k��^��!W�����'�L
�Ā���8A9�o�W�3v�V�}S��7n�+
�T]�r��b�;�+�!|����)oٷ���/A�Q�P��5V'ᜳ�;2�]��+�OM�l�`��@�3%"DGq�t��.��}��gH[�^�3�4�nl�׫�kL���K�ދ(��o��ek� ��#�$�Tk��J�nn$��"{�+Uv}|2�m�-f�A�o�'��8��KU�	Uqz	��j��bN�ET��9�0ܞR�[����i���;Řc��	�(w�)��]�$c�Jɮ��I0������Nq��g��7����2R��!|;L���]��,>���?�'j��"�#����C	���ٛ(��s(gt>˄��8��^͊�s���_$�A:���oOњ@�@�1B���фN?��#���p��;im(�Qn�S�r`������x�����G�ן
~��
	]	t�deoխD.*�I	F�z���.,`t�_4&�����x��ڞ�����dy��q,��[׃���1�c��e`��[k��< �{�T��)�'&������� �D���Ժ���&�d�J�QY�d�t���}�	����?���K��:G+4QF;୆�[��B��"I0�ٗ����~�:h���xN�ζc~�F�F��?$qr����6+�?�U�J�����F���\Q�F3�02�H��Q�^�1���^[�����^�^�}W5��l��������S���T�j�K�ܧ5��?΀����p%^���ل6Ψ4�ן�p��M }�R?M���x'l��f5j��X�iT���B�#����~�85�����[p����~��hɱ2cF9��п�D�цW'Y.�)�J�,�๼�-x�������5����oxwZ��ݒY�{����k��O�$����$ ���f�u�Ժ�"L�XG��x�C`ETW.���۫��$��0v�&:������.׳��7�bB_���	 ǽ�;�3 �;��	��[Pvy'����RZ*Ȩ_,N�3¬��(l�.�&U����n����u������0z���2���.�x�4͚����w �v�U��V���.�N:��Gz�2]{�},�t�1$e�K^�"�p��g<�G����3e �	JaoҼ:�V����U���?uă��G{@O'�aw���-^nד��I�}C|���;���yc�#�����5��l58�$jp��Ge�y��z���y7�x�[|���ȉP�S��zSs��KDI�L[�J��Gw�F�����j>h�́=�O%�3�c��w9�_�^�ȶj���=��K�-~
�t<�a4�C�=��H�[��k>Zǃ�a�e�G�d՚��p%��pO�|i�σ�˸t�ƿ#V7���y�^~5}���.
T��<��Ā�
c1rS(.�[�	�\s������8� 4�x�Мs��RJ�l4��	�1�a�g�_�7uT�����
���I �r����CT�z��n�o4f�L��3���n��� �~|>D�|��8�;i%�E�3*����-�D����ʢ���c���$��H<�\Xgdߔ+p,J��l'���1�Y����0�̝%R��3VR�53D`tY'���ȭ �Ph��1�ݼ>�gf�X=X{ۙ>;�4�؟��z���7s�m�ZV�B�M�e���>���#�tdl$̉�Se(�Ga�}��&�G��"�OAv�n4hf �
�L�-E�- ��H�/��I�$���V���*�Q���� ]�a"_�q3�I7�3w�Y ;�P{��� �4m�iQ8�.EF����;�����XZ՜�w~�j��\N�VN��9g��*����&�ս!2uΑ��"���Ҥf{aW{"��z����&��\��TOw$.Y,Cz�"����#�#p�xGq�
^Z��Gz��_\���.�����ll@3s�+8��[=�l>v�Oجm0߀����楼�8D��4{����+�L`7��t%���0 ��uk�TR:]q8��{�8*��R��n&V�4��c�P]4�Dd���򱂃�%�b�����8����@�!n��Kbc͇@V�O���YI|����=t��>+�<2w�)
�ƽ@~��.䤼]P�FЍHu��6�Q��� h��B;�n�(f>�C�Mw51uߟr��~��K���e~f�7R�,��ϼ���z����(Vrkr���l�N��.�xZ#^� �:��^i�=-PU��Y_+!N�Kk��v}�RI�r���/��޹L$JgExD����/U(�����f�Imf1=�݉�r��Q���
e�hu�Xo�+��g<va���ծ��~J`W_�� �Ux�)�yY�f��?݃��W�(�_K� =H�Q�j�x�;=�b��E�:�:Y:�w$5{6�ƌ���=ɴ��9��^�E��c��iSo��� �r�&��D+Ś���w�Vm�ݫ�%��R��Sp��Ҩ�>l�z&�	�ܲH�m�IVҔt�	��k�Jc3�p�j�F�^��Hjx����O'���Xq�}�9�+�sU]���3/���V���
�c� Ք���`!�&A��tio�/Q1V0^�~t��\�Z)�j��Q�a�Y��~�����e��Zr0�J,4n"@[Woy!��z�,grO�A�u.�I�O ����"�,$"%>���?ڧ��-��Si�����������Q�+0� 	y�9h��Uw�"CPڵ�d�)F���*j��W�}t���B�L�U�1�Ȭ!c���9�s��>� `��D*\�K%�?��g(T�+j�p��)����B�$��7��+�����l�r'P\2`�;�����'5�+�!��WG�ҏ�Rlz�G�|�8�J���f�����9�H/s�i�Ȝ����R�s�T?c*���2��p�5��lt�94��b��0V0��f���p�}�)ҭ;���W�U7Ğ��V���w�G�M��GQ!��&2�'���o�S�&q���}�c���B�=7<�����'1��]��8�y����!d5S�C�(�����Z�9�߶�1NLr��u֡	��qt��^�r8d�CrF&�C+�ga��)|T�֣&Gͮ�YVkGb,���n��ﱌ�p�W�����T���~a[E/���1���m=�J�௣� �BQF�<�FFi�Tt��)�]�H��"�6�`ݽ� "���ׇ%m!wg�X#r.)��B\a��xg�s�
���r��nn�&uxBS�B%�|e8dOdx�#Ҏ�M?�"�Nn�!�줢��߻�ͼC�Pز�z�}3{��WH��@�}Ѝ�n�
U�4Wz_�'R�Q��F�H�)pWf�P�q¤V���V��5���$=��|T��k��Mأlv	.���T��\��Y��m<�J3���B�.��/,�����8LQ�b)�mM{�������?���y�(Ms�!Z)o�����r��@��#)8���^>7,S�Lv�%M����lϧ�L��QbWC'Ϥi��R'[����r��eʗ�T�䔖Qۚ]�����f]�����un7�AI�f,Ja���Oh������ōyNZ�E�����Sj�{��g�hS1��Eɠ���/���V�"����,��6"��k(1��A#�� ��\x8��f�1�}�P�s�6c �����]3�ZS�m ��֔%Rc-�ds���k,�*x�:�Y�i�e������WoD�!y �VëX�1�X�X8i�Y'��2�[`��v�Iߑᯱ���Y���/��X�j�ݖ�,ŵt4�(Fz��$��(I�� M���x����]UG3e6V|!]�L^�H�$%�*UEG�PZ�ɑB�X*9�K��)A����/��quD805�\�Z	?&�d�:�Q�O �Q�&|<]����3haI㸡Pp�8>]����P�c�)��3��PW�2#���W!f��0��G��j���ɮ �@�e�`��S����y-J�נBG���Y�2Y���X���&��-%�o��>&9dH8��_�3�y�d��y��nd
d���~4$j� ���Ѧ+��We�Ř�I��P�����d.}����Ŕ~����F2�^4�ʛ�_���@b>�TY9�y�.��ta��\8ĺ��B��.�0�I����df���$'��2�v���I�P|Fx}� �/#����0o2P�&�NBT�^��M���B�6,�3*w��<�6��?E�=qa�pQ�Ŕ/�<�~�2d]�#���P�'��r^$�9����c^O��޽�~q���EP��M~L;q���*Z�hG6��E��%J�4h��O򚷚�?Ƿ?�&�e��d��Q��@�����h��O8�Bb�Y��3
��AZe»�R}��67�aP�L?��8��m@��BK^�'�Ou�3�?S��J�+���5y7�]s$\8)�R����V����\����~��i�,��2ύ#2��JM�+��E9��_�놙(�ƭס`ؗR�-OM`w��I���2tZI<��
5��rT�U�6I�ԇzubA����]R\H$�7Q�<������0&zz�3���Ա7�ݟ�Tv�nZΕ������? �~$��Iy�3T�pT�GC-�t��7Q��ἃ<9 ��pw������	�&RM3沚S�Ӝk�Z<9�\s�$;u�`~Iќ�`':�_f�>iyD�<�H~d��]g�������r�6���b����}���2�x�z	*���������Ib-*m6��� 1;R�B��"	<�AK�����8���=����F0�Y��Z�Ο7�Yk�\>�y��P���B���r��~�[&e�(���`�J��W����=a�3�#G�Æ}>�(�}���X�1:���1��ۚ��4�AE>g�1�(�
GQ�v7kĖˡ�I�x�M�#�>��\�IFS�>7b�=��	�J�����d�v��)5B��J�a�F��x2�� ��<���m=�<��W��Y�%������D�	'}A�³:�?�ǃ��2e��EL\�z�X��[q%S�VQ_n2�K~�l��!oJ��C�"L'�'��Ǎ��9�k*���P���j��/#�2hm{_�A��+9Vc�բ��ZRf�Ɖ�n
�^�h!񆈩�����[�0�q  �.��\ �2v����8H6�ND���D��K��p}�D^ h��Lnڂ|ш~;����Ȧ�&}���r��8(zm(�`� ���?�[&��8b'�@���[A��3�р�d�)�������sE�i��/����,�O����H��3X-�X%��VF��v������"���Q�%�{�t��/(��)���Ϲ�o�x��՟�If%JRʗQ��?��i+Į(8��*����X+8�كx�&/�W�w���4��[�_W%v�a�K]vf�!���P M7�+dz`��hR������e^`uU��uȍȠ�O-�ֿ��m]�]���Ӎ�a7��g�f|��1-�$[��m���Sn� w[V�iޭ�wE {��XaLu����H�����d6�% ���&Z�z�XC���H�9�^<��5T�` �2�m�6�Y�i����N)�u�XP� �ȫ�+�g�ҷ�SG2܌�'�@���8fK �^r�vY���\lX��-�A���:����Uy4���}�Yd��GAG-�z"[`����aH7Z��=Y�拇	o*���d����b������Y2G_��{�vN&�mxc�l����ݦE�E/)�' C��?�D�\��;L�h�yLu1P����X$�א�i����Ou9�#������)�|SB��Z�D�PQ|���P(�Q���`��1�U�E�0�y�a�9��,k���H���pt��������9�e��EY�D���#�P<�/�|�A��f��t%��뫳�öɻ�Y�	q�x�v�ls���FT�G�
0!�pCk���H��b9�5*�i6)�w˩
̟74�o]T��l[��y��p�l�7G�2���������w�������B	S���y���}-����]�Lq7�\��䀨���)�R�Tg""آI��_�<���`v�l<��a�Kx�]�=�D����}`���D<��#/���K��I��l��ߞ���,Zo�����s�џg��k���e��7jM�ak��z��V��~�.��Z8# <�:�&�
�#����;F�!2�x��oae�8v"��o�c���}�wcU�ӟ9ME��-��И��/:�� ���B�6����	l!�R�>Ϋ�o���ݯ-S O�H�b?�0IW��D�ԩ��57�qn8��\���0��,���W����	m�˖ēva�e�Eq"Iw �hm��l|]{���t�5���W0u�S���<�먧oR�<-�U 	�J���'Y
��� :Qp�nB�cYq���!	�G
МM�"Fv�4I�Z��ޮܿB�g�&��%�%� ��"j�=	��n�H��;�`OJ���;��Z�K5��坃�c�h�J�z��H؃��l4ꯌ�+��hj��RMhމ�:���`���v��ՑS	ﰉ1���b��?Gq�"��D���?�P|^O��05�d���6���А	��{����a��Ӭ�O~m�K����aUE"����Ϙuh�.u��TU\L�I*Q��v�oc>M������j���t��� ���h��p��b.T�����tl� ��4M�V�A�*����O]���->6�r���l)	;��p�UA�X���y�'v�b$�����h�w�xu��x;u�*��ަZ�7������	��-I12G7�A���ٟ*���e غ����[~�#�Ir�u��gt�`��Y�.����bo��%�8�r��� x�7�!
�1��s��&,C?�a�E�BW��]]��-�_���ť���n;A�*r+�s�˚E�T�,�b�������y!]?4�'%�-�?ҁI��N�,t�I������G�T�
�H�|�>Yy ��S��+S�E0ǻq��j��~}cw�7��)�و�6E�����.f،��Z�.szN|���Je}4~��o!2��/��wd��¿���@�%�:��|��mbD�ɤƪ�V��x�q]��Q`�]d�oDa�Ok PA��-r�au��Z�6l�"�x�\x^sC��I�Ѡ�Λ��&�+��y�@�ϖ�\�(���[�UX9Z$V��f�?�ǯ�lE r5��@{��J�����������R��Ok�_�'��^vB�f4�����:Z��!;���""?�q�mlg��z�� Mo���7�}"�F�XO���#�͈Zso���3�k՘�i��F)�+�m�ʬ��ܑ�l�MCl,���Ń"z�4G-	���V��m��Ț��{:��BK�qL	Z�]�R>Eg�Y�E&�$l%��غ뫄#��n?�%w���C�&$�]��hM��x]�P�ސ�l��+��~�T9y�k��*Eu�K,�<H����AL	%�� &\���g-LB.�[�n塲 h�#�����s�{�e��u��P�6 Y=o_�(���&������?��U�p!�vn��F���E� µ�_�������3�*x<C�Z0�c�xV0�����&�0�O���v���\��ւ�gr�蓵ԁ�Jp�(��~�)bCL.t֍�	=�e�x�	���.+�dd�~Zo@t���s�jt��k�Ȩ��qKEPGbU"t�Ǝ#\�J�oU��R�=�e�Xj�&p�cD�Y���@�lÀS^��d��]�˭!]�d�2�l�O/ !,�p76\S7�E2O-ґ+]0��D3��]�Ƴ�>����?'�8F0\18!7��&��g뚪9!�n����yI���������.3�HT
!L����\�ͺ}+��.X�8ggJճA~�Ez.9]T>}�^o����@!����j�a�c�`Fiy�O�<hO|��$ۋ�Xӳ9+zd�-�^ߢۮ�:�i'��I���z���º�fo#�X?�I���z�H�L���Lx�zE�#��oJH�aGl��R&��: :(�n�D�P�TQz��H��Q��y\�~FP�/b� '��h�6H5fH�>���~���v����"���Zv
��#S�,8�~��<Ѯ�I7�&vڶ���AJf�l]���o�@�rf�p
���貖!�A���ЫMMd�hY�} d�%ǅ��_�ЄH�yd3n��������(�6B�L�(I�@�.��ü8�[3�i�U��Ϯ���Z���Ej`߂��kI���^2�?����dK���n	T�[���Op0	�Is��Z �s{Ƶh:[�S�٬���(��K��c��m�^��D����>�P���)���J�=����=ţ�]����W��Ƕ�M¤��h�&�[{��m�i�v!E%l�12�6��?E$Ғ\���ڶ���9Q�B@�]rt�+���4?�%��!-��;@!�>�l���b?�/Qw����[��P�N��"�
���ҩ7��so5J�Q�����SyJ�>�� v�N��;��5n� Lu 3������~	�!��t�\o*37�[p�W$�"'�/Ϸ�Կ��&z��O�h���8'F�s��<�0�C�s	�@>�}��	Ǩ``�U�喤��վ�l
z{���5��),$���K2�S���I�Y��B�2A�<��@7��$-l��=(�(���ҥ��y��#-��#%$��E�Q4��� .�A\��|C�Ě6��n���Ic�Y��
�/(��	;� ��U�nj��z� ��6JExh�5��[u��٪A0�ަ_��_ί������A�X���N'eq��_ϛ��b>�_ݿ%b��w���`{�z���c�Z�#�:��M�9x��j��Du�E[���S��j_� �g+) E��2�I�͙���/�ʗ�w�_U���'>9�Do<�u)�@Uڽl�,)�åq5����v��^;���A̍/�W.��"X���u��.[|� ���>�C�u.=�������o��􁝮��xǠ�-z�$ۗ���U�Ʉ�9pH�^"����?&�Fld�\��߹�Q�V�0�*.��S�j7�D�M�yȔ�������?�ϓ��
:,���G#EA��d��`w��C_�����;�jqU�v�G��A�m �{ 3�1V���O�TN�^��`*�2JB�E�ہj�LM�� �����+∣ܠ�W���_ogWv����
�gF<�%uh��3P{uY.����d�m-N4�M���)I8o�V�?�1^��h��z�d�%�0�C^[3꞊���z
&�br�����cz�����6��>.yW��z���Ws5O��f /�?��X�v\dNϏrg�S�VS/���y����{sU�<f�~#Sp��r;͙l�(���|�К�E,4�/���o�t%d�\�zd^Gd|�����a�iG�q�)kx&�9�j�Z$Oy�� �(Yx�F�tCP����E1�~��.��}�}��"�@x�n�R�:X���,T(dn�`���ґop,���}���,�A��@�d�Ǩy3ZJe��-o�o*2�]���^T��u�7(P^6�{��W�k�@s�i���uJW�8|����N-���䞽�nj��K��Gv��5�����|r+F���<M�^�4�$�fk���m�M����v��.s��{��ާ�KÄg�~E�W�k�jc�d>j@X!����`����ױ�t��}�bS��j�sL|�-���ۃ,�{�%:;I-Hkwl�8"�� w��¸������˔���/��2�w5 ,~�a������7��e ���TV4�:���H��C9�PM:��ER�{!����]���״񜌢�TO$����q=����uپ�:&�$�s�id;W�������Tq�og&;��}��8���b�⇦�KET�699��>b�=�Z�F���zq��B/M���.��W-7Wx���a�a�����������[�<�ۑ]΋Od�V��|56	k;����K��t2Q1�a�n�OD)��q��lOu.ѵ�z�ϫgc����$X����ۍ��y�/���F���
��W3��a)pr�`ڇ���hY��0����)���rq��g���@�n�3	j�にO�Z��П�{矼r|�)7����xT3�Q�B��mgd��k۷L�e�/�U��,�fcˡ��������>"P���(�-dMw3�w~�[��d�T��1�8�(�2Q`�8ա���M�,kp)�5.�!�b��؃��W]�f��K�-%���r��<��fF5���U�yc�=S�ܚ�N���fZ"3L#�r��s���T�0�������3��BE7�-F�(��|[��\���}0��`
�n�]/��������Ł��@g�nG��8'a"�(8�� Ml�`�Z	�b8��l˚�t-�0�x^�yV�)��9^J�.K�^�bxx�G� ]ڡǝ�Aȧ ���3<a��'���A�5���9U5/������4��0+m�Y��]�X0:��[�׮A��'��7Ӻ�'���V��:�B_�3_�qA �)��1�и�Y1��C��!T!0����k��xl�¤�q�Y���VY�nGHK����ި�kBቲs�6*��X�x6��ϑH�N	�R��q����]��L�v�\��n� m���,�������9Y�N�-b�l�m�B��Z�R#�d�%봲�**�)%���cWI("�KLn��.����
I.���q�f���  
��)�"u��R�v�����y��w5�m1*oh�W����pfwuM�I���,y%��D ��VO�����}7#w�e�'r?�k��4�1u�C��Ċ���`�=9�u#�� S9FLy/�x���t�ݪ�7������Jp����i�wʷgk}\�'��0�T^.��$�qM?0��)Mz9���j
�#�u+��[`	��s��K�.?��8��� M`@���f��:�����/�"��컢Ri>i����˛4!)���
g~�~��Bi�u��~������c�$g�(k9-<�'"�ç���y��I��)��\�υ�4����l0�{��߳�>�ƅ�����J�*[�87x��I����쫳�e��X�5A�_m텬GZȴ���k�x,����]n�����d�i5�$����_%�uC��@�\��D~ov@lM���/%:q�D�I�@�L(I
����;�O [��aІ�:D�l���;���;�<s�K����b�
�g�-8i�U���0��-je8�sK2�:�ťz�I���d�7�G�ʒ窑^�CQG�L=�jDd��)�1���H[���6<�'#ĉ!��5�MJ�c_^�5�u�_�`�^����A������l�Φ.�Μ��h'��^�m�g⽴J^�A,���>|",{��Y])?f�� 
�~�/)��v0�A��
�q�R^�� ��6MWxdg�K��4�p�O���aR9Z��@ה�u/^.�_(8�J�MK�1�t���������QXʰ�l ���ʘ����MhV:5=��!\�:���
�ߋfr�}�X־С���9�]r����9�y!���m<c�;oJ�8��2���`�#���аe�%�q��pP@hI/���'ӸΗ�I_�*���Ȩ�(fGx0B�=�7���fbV�Nr�!
��v?�4����=��-����B~oǶ���`v��YeO���2���HBV>N��gm��$K�g� ^��\����id�2��� 	�捂��o�������$Ip~uHW��2B�!�
O�>���\�z�4�Q 5�L�[?�<����y�<��M��k�#zA�M�\�NA䚍>����$�����n������>
���L0��1��N߭a#�eɷ+�i���zS�E��x�N�}�²��m~�BG0/U�x�4/���^�saB��$�䌨4����%�{PN��)�>���y��B 8���/BY�vF edr��V��_���s�y�z}����>��Aw�.T�#����.bNa��u���z���|��-64 Xx�0Y3:A�i��m�7-^�4w�:_r젱����HJIX�/El�0�RݸC�T'����w3��lT��Y�Vȇͫy���`�Ji��T��ZF49�aV*`�o��x��Z!C,��Ҍ���o���X�K�#����N�gE�>��E���)Rwp�E����`��ҡ!��&�'J-?����E��Kx-�����h}4�*%�ԭ�&�:?`������Գ��2��bP����	����v7$�lS�wAz�1U��)>�����G�#_2C͓P}{߽x�~8���o�!� ]+,�?N�(gL9�Ȣ7<5f�^8H*פǘL�e������
	�B����8�$�U1~�9��x��@Y����M�4�U8'%G}�e��zJ���D����{#ΐ���Y�Jy �t\�{��g2!ә�Ά�_,T��֑~����\��t	S�j1)�ݬCbҧ9�7�I�3:6��͔�K�7=�M�j7!=/p�7j�wP�YN�Ԉt ���)$>� 
�L�kD�i�u�]�_S�ǝ���V���bZB�i�R���K�����
�E9�%�;n���h�25� r��c� �a	s���J�hḽ;��9�ܔ�B�����9�F����!_K�,�S���W^H,�2����ռ�C��P�
�4��i�Gm]��h�L+5qS�{r4QL�c�
i�f��6�*OI���Br��O �T9��"M^�,@�7�ӽ���<�b����a�S�n��2��{
 V�,�
�;D����-#�j����w蹌�O�'z��o����%.T�6�!]�H����{3W��58�?"�a�ѸxԥK?��#��7d&����PP?��5���r�|d�zG�i�.=��3g�}kx�R��o O��r��"ѻ�s���X�:\XL�M�m�h�#�u�/Mb3	�F���.KJ�L��"��/���j�F�U��6X8� ��+�`�%G��. �-����Cj6# Σ%j7���8
)$���|uF�SȎ��.d�Hoc�aO^QKѪ�ьƂ�� -72��}�舵���Q:_�y�[����<cDo���K3�~�L�����WIkb����x�^�hDN���<�q�������vs�`B���y�
�+���Ȯ�{v9P��L�(vs�G�Җ�<��|�Obإ�?�C�F���;2��]��R�d$71aڌ7+(WD���4�?mt�
`��îAdWe_��]����8���3-�k1'͘�W�Rsp`��Ơ���au�^��|/��O<������Ԩ�5ר1�*�c~��Hk��]�TEA���02^MNw�/��UB+e*^�D��_�k|����6��Y3�2��360-�����b2Y|H���JS�| �����D��x��ޱ�C*��΂C�����n4�l}����N��"�>���-��+��(_�ӡ��/�
r����f�RNmV�G����.���t����XaH������:8b�G���16��d�Ǧ{I5F���t]�ϛ�ݱ��P�_R ̠���9���_+}WB�2<sy�� �y��N%�Vߔ�Y_�Fl�	��3_'M5D������	�����s�A�߳�W�V���Ew��gJʁ�>�t������*�↿q����
�u*�l�1���@�̓f�:��
��:6N�����c�m��(SVÕlD}��G9�����"p/m$4����.��&�$�+�'��ntU;N�8���V}��Bg~��Vռs���7|h��B��W Z/��x��@��7�5^��3�<d8`�
zU]4��n�wtCn���� ŘWK���#�+ny<�o^*yP�^G;�[���D�T�c2W�nڞ� a�Hч����e��
1�@�4f�E�����i�6����?�cMG���.����t��ӂ
߳��ȗq:8x�M +��*��V�ƝѦKq^P$��ϴ�w3��j]e�焳�G�?DИ)Y�Ϋ�8Yo+�p�j��y�F�sbe��/��Sz��:�k��n���@��Y�z��e-�H��b��q�O0à=п�Y_>���L;u$��Y|�,m�9�+x(�&��?�s�^W'���,uwU=1��S���[���J�p*X\�ط��ώaN�o3��E�܇�Iq6�ɂi#0+ϗ�A�`m�B�p���m͘H!Jպ����%�����Z0OFb!(ל)��s�9�a�f��8~Y�#��K+�>�aM�������>{���w��ۅԻ���^��A�8��0.A� ��d�\��OD�U�/��R�Gzj��u+q�{��/b���	o>ǒo�M��u��抪\_O�z��������	��c_%%�q��_�!��6���_P��6g�T��c��T�P0
ي���2L�	��]������:X��O���
��[_5H\^`N7�:�k�-��`�?�Mt�xՄ�=����A@IںZ�ۆ�0�~=	 b~W#�+����R�6J��#�vB��M�@>Ux1��2t�`��*����Ԃ�vÃ�ٳ:�ċ8~���9=�\��_���ܧ_5C@Zp�2`��N˅���l�w��N�f`�����]y]bH���m4�T|�8�:��̇�����8�3����D�>�H��=45���F�����`nf�	0�{��o�G�]B��=:��r��_Dw�����r�����v���^R���G-D4	��W�D�����((a�\��.�F�}�#�'Nc��8Zn����)�;w�5�3F^(���L�w���Ƹ�lv&�繙Z�]�ї���YS��Yx
��>%�Œ��� �N=	:�oa�s�zM���<���z��,~�X۹��(� �FN?,C�J�{zEot,(<��ֲ(fR�Fy����B�a�W�H�TԛW���{r��!�o	>-�[.���W�6>̀�(%�G2͌2}�cM<�@�4e}�l4�O�Ծ���^�C�`���s�W��A#H����#�0�`ٳox��q����t�,0��Z�Q��(����X��W�w�5n
�eT����1�W��c��u��������9�P�[_�6���E�M���mu�����Bvg e-���vZ珸�8��Ar��;��]�I5�i��>+� �l��d� 9vv�Rq�.�QW,�L�U��v$�����4>��L��K(�z�$��!硝F���ㄲ>��̣�>S��eMО룴1ŝɔ�6P�e���x�{c}�>��,|�ՀoA^��5��6N��Hhv@z_���MCe�%:}��Cuh�qk�R9�hmG�r��CCF�w�pb�{���������q�GE_
�6��������5N�lھ�=���i-��t�����Y�Я��<"�?u��+01����Ig�LS7�ұ調IYg8'��?{���'ئ�E�B��o��f�9ѧ`#J"F�-����S>(v�kXT��J� b�/��+]���Nc<�R�߇!���)>�tд���6�'�OCd�V8�e�Cڢ��x3�Z�j���#+j�G~�lbN�ehp��滚?�='SP����x-��i(���k�e�R���J���W[���
�� }��ײ��W�DNkoU��	�:�ĸ�C���+�I�Ġ�A�Z=�a�����/�5��|����oXcus���d�59 ��ʼ'�j��n� �Y��#�.���g\���0�jE��F+��	VH�V�����0����*d�U�sIsT�T��4�o�o6��u[[Z�"�Ӫ�n�d|a�
mmĨ�r�A�+�e:���r��v��r<ي�ٓ��r���	۹�Xu�3�"ɦ^)�=K�_���74���>�e8D�x:0#��r�Z����h�@��_�On���d_�U�z�}��'`�7��*��w`wĀ���|ǟ�.��oS���I<�P5<
��x*��4t�G�!!�	���Gl��u�N��1�4x��7D�m�s���3���+t��Ng�'���,�-�ﺦ�}
�D��U������rQD|���F�B�_��,��>�yݵm疴/�RY�2��.����b�2�1�L�ZvM} l�-T���P�ܽ�O�Z��,䑢�g� ��Nr�*�s.ɕP�8[G%V5�8��*jZf}�b�Nh}��`�\bW��fތ�\�g��G������s�L���+#:�t���P�w�Sz}�\39��ޠ�ݡ�M� �#9i��+�:�M�tt�?�=Ζ��[������¦w��������_� R�9֯����,nL�3��{�f:�F$4lo�y�h�zJ��1��O7+f��ʱa
��E�K)]�x��?�����������J�?�
lc4�����#�y�d�ͺi��*�ܻ�n<e��c�k��n�ʧ���Ŀ_+W&/0 <������v�yШ�Y�#^�W��l}�'˙��(|�,�����n�ػ�qi�����X��~`k��	kI�8�M-C7����}Ơ!;)GK�D��I_.����1���/>���a>�dG*�u��i!�9gS��9����7��E�G�_̄!wʭ}�W3��nE�v�Ψr2I��E��:�2��x�.���\�D�?�� �p�[h��=���u��%�s^q��.�
���u�1�2�O�y塧Ǖ��K� }i��GN������
�M���������I�1���(*���þC��("\�x�ǩU���D�{��x�ўX'���{
3�L�i0wH�^� �qS�#Q4����C(<�A��t�����8�s"+ld0S7��/cl�^0o&�^j�I`��� }w�Q����g����H����G+Gt��i{�ť�A.Uxd~g����,Zڛ�Y�X��lU}�z��%jD(�:[N�۳��߈U���#N�x���2$���������jN��@h��.�)7�i�nv(��{C�e��J�@��h(��t�r��i44��Kvh�ٯ�
�#(sݑ\��*��A��Bȋ�͗�J_����@��L�/��߹oRQ&�շ��
��d�h� BS/����U�D��n��|O�?xD��T��=�/�w�;d:�*k����?���B]���ninI�H.$	�W�}-l܉���y�b�)va�?��8����;p�|Jힶn��هF��ѵ�7��ty����`թZ����	����o�=/�<I\�����v"![��cB��m�saM�����.�K+_7��&*����cl�[]�V�C۴�6e���4��~����9Z��\]Y���DC�ߗ#���)§O����k���u���[�.+|�\�?�I-d�֏��\h����㞮T���/��ěQn�����#i�{�dӨ3�2�9����:�ɲ#���mV�В��`����4�� G�f�"?^�[�/4�xk�=�/�>�I<7M+�ϡ��*��َ��@�ߛ�~@\��g���d.aa�|`_S�/�����k��H����p����_��T�[T������'�_g])���WOº�p ʮ{g�`0B�����EP�)�W����I%�&��*��y��a��G��/9\U�i�L�ί@ �]�Job_~g$H?Dt�� T �G,���
�8��^x�Ғ;����2%���Y�|���,���zBhOj��'\����x���T�D�D4Xo���dvg�:3UP�S�צ�T�x��)
q����d��n�D�>nL�c\i�����ܑ�>��:�Ճ�c�@�3��.��_u��lέI�	�<M)_�)n|�����V	_o�ߞ���Jh�l��.�,�e����l]��_����}W�T�\�m2>��U����.[�5wb����T���\�vX�� aħn;U^�0�`$6�kDP��犒��F%�?r��;�⇺S�52g}�\<�fS�?$Xl�K����f�|�\Z���5OJP��0���ٿ(!u�ð:s]���a�w�5d�F�^"����9e�U,����&`ޅ+A��Ԓ�����Żh��1	��=��#K���dˊxL���,���T�G`l��s�/#F
��Ӥe��:�0�P./���⡪�yS׆����n�Y�V�Q|�V� ��q�u�qQY��D����Ç�nk[��>�	�^��	lPv�J�爜RQ��FO�O�G�w�8R,md%ݱ>�9����Lg�lP����x�;�i�K��P��/��By���R1o��5�� &����'csPM�*Ku���sy��:S�5�����|ݦ௒@�e>i�9c'<���$�J�ئ�.q�����3htC;m�9|'��B *�I����;�և��&��-h�q�T�_��h�Ad�z7�L��t9���s��LiM<��h��66�����C��I%F���Λ�>Pb��4��Y��KnK�_�8�h
��އdNk���[!Yf�͡=�������e�9��j7=I�Ak��r�o)8�)� �,��w!�� v-��׎I�˩���Gb���+J0�k�Ab��)U�aT%�;W)�����B��]T��_2�a�x$���\0��h��m�H�C��i>��]��y�v��_Pfa[���hH�*@��n��_���9g�{#��k@k�$�-!�b�t� 	�zC�ܺ��g�І?V�:�D���.:�3�4�lؔ�-4ǘ�SٓX���W|��V�G�x_I4`�[���ĪKyăT�
�|�G �a�#i����Tp�o��*����q���ܚ� �Z�<��,�J7�G�K��HW�;�>-�����(j�S��FGl~�����щ�ݍ�Ϯ� Q�\]� o�����8S�.��,u(�>��'	�vi�@J%��ps��V��ݜ������d��9�����
��n'L="���(O��o�k�8uY�<y',�i����R`��fϧ�f�*0���ے<�)�$�+XZ�@]���}��9y��ܺ��L��(�޾�]�J���_���B�j�b��԰���k�����uI�m���F�`����L���Q&؍q}5A��y���C��?f�|K�����}��ʢY��n�Kn�Ė�̕��A������t%꺈<��f�`���6F���2�����4 �>jY$��l��/��ś&Z\g'2�$X���Z�����.��6��uiPy2���QDU�ʲF�	$��Jd!��ϧ�~�P��8Vh@/����dÉ��BS;��i���r�C�;a*JV{��Z`aQ���p#6ei��eJ�h�O���R��"�L��c7��'���F�C�f����vhj��`�4J�!�)����:S4�'ϛ���ц�ɾ+�t*��k�D\��1��¶�����a��a���K铐Bo�HU�Kh�&7��-T�E�b��Aೱ_� h	7��	XTҐ��l}N�U��:kvnF�.C�Y��Ħ��N\U�*9aɟ�ˏ]Em(��2�bE ���Q_"�C�r���6i�T�L;�ɫ�O-*�B�ᅁ2>�HP���HnPN��Av��������#�.pT΃����j�2U|�d/m���݅f�2+̬r>����H�}?%Y��
3:Ⱦ��eK�23�P��Ӆ��}T	��$�u9.>Wb`C�H�R�IòoY�P
Y9T�K�f����7��_���ڬ����$7
t�)�󺱐��ȼ|NW~��� :�����Ht9��Gʫ��RPi��	�0����9��!�h`���cV�$�%�_͑ܮ�9�!�{�_	�od���,�쒅�@S"�%�� ��o:'�u�4)Yӓ����S&�5�@y�v����`�]Fj���>�Q�#�ƙrAjA��!���G1�(	�@Kh��\'
����"�Y3�� Ql��Q�A�x@n�H�o*�2В���/�?J�����M�˼pXL�׫K9�ڢ�9�l�u���Q�#u){�N����|)v�/��_��j�T]t�ZZ�w�0M��y˧]P z�`�EVg��Ƨ@g5�>�W�h�� ��٬n� ��s>R��jJDGk��b1L���f0���͚�ҋQ���d�UÞ@ZAbZ�n�Kykj� �n�۔/���׷5s�x��r��kO��,��a�h�Xx��� /��OtZ;	�ֵ�4������S��kS��u���wZ�z��l���Ǔω!��z��Q�:j�U�A0lj��r�3�� �1MD� �.[C'��3���-a$FR���-eZ�.4��$'ը"��(1��ľ�<��x�WQ[V��cX��Z�T��_ 	&��?�T�O<�P�u.�=��$[YS(qE�j߃x��F��6� ҏ�N��l=����I���B�љ5�k���(�R�-s�\!3�O�N�Q�����79�#�����Z|q��C#�����g��?�ᐞm�Iͤ�Jl#��t%�L�y�^��{H�Ko��K���Z�5�ܲn�E�j�O7��R��<,Jp���_i���UBs������Y��d�!"$b�1�}�)Y�Yw����3�1n-`
�U�ՇL�s�1���߃� �e��0��C�V�e��ؐa	1^�x�h�S5�qd��&-%��g��F���LR�ըrt��S0`1^9��ܳ�*z���Vi�Y`�^D�+� ����	R�ɼdh�#K��ٮ���������)�\��q�jE�3�z&D�5�z5s�,��c�B
�
��ě�2�L�9������~�j�S��E@-0�O��a�L+,�+�A@��!��fF�~�ټ]�{H:t����UpJ=����S���
�q��,�!��,��n���E�;CG�U�Y0��!���\��b�f����a�um+Af���1v!>��E��~��=P<�H�t�)��;̄�^��:�$� ?t�%�W�ڞ�p�{�=>���B�Φo����1��֕.B,��И��[�Q;�(,a>���?L�T�΃"������/�~�X�
�7T= `_'S2���k'��.��E-|o�f��g��B�oc�#TU?�Z�����`��mE}- ��`��W�Pci�z4�G��d�9��������G\��F��h��/�
gN~	�]�Igq�XGCC``���?~�y��}���
ܪ�J����F�̥�N���&�t@w�9g�S��Q����g.���*,@���VcҕP�z���Ln�����&�ϼԿ���gD�g�!�%r���L�$۷@�'�V�����~waD�yK��Hȹ?���� 朵f9�kv�+Z1�$0}����(��j���s͇�귝��SzhLT���]�"��p������/\s���lD�U|�0��<I�ɧ����'��;,��C�f��?J��E1c�3}���<%۶��F6{ �ғ��m�·KI������t���G�!#u(o��o!��eڹ,n����4�}C��c�xg����G!�=�"z��Q�`���&���#�T@�˫.ZT������$��a#�u���YDii|�!��öt�x�Y��*utHRn�{�T�p,6�[A�7S2ȧ�9�g�HB�T{���Q�*W�`�
Q�-�P�xmh����8��	��qŷ��>��;w���$6Í4~��C��K Ӏu���bN`�|uN�N��XX�l(W�� ���p�l�4W<�m�H����e��=8���J�s|��9+CAVE��5�����o�^�|76�㓣�N��ь�
�T?P�i��I�px��#�h�>������p��'s�a��Fp1��G��A�`��Um��(�����BI0σ�1^Q���;���r
[q�f�3�ɠ�W$���ݺnv��/�Rn�3�U�7]D����:��$Ƽ�
l_��F�\ٖ�^����TB��[7f�Ǻާ4C<��#�=Nk�#�����2��aW��铊!�Я�Ȋ��w��mwP�y��2@���ϑ�(��>�X�=�	%����R��%o�����J��Ƃ�B���[��Qx�M���[M�AR"\��j��@3���jh;*e+�%�R;4���Di��=J_&�dD�*��D$�N�:��Y��#"Z���M��}̝��F4JB�ҘaGT�>>TH�ٹ������B�#ؒ-'�ZRC|B����kg@s��It���H��ZO\��"�%)I��u~7���ru�9��t6-����nY�C����a4�?�P�\9��he��#��«��9����y���a���_��?O��1զ�r�άF7�3��t[�4@�،5�����gz,-.B�d�W�P��:*i����U�^���m�|dr3���|��o�}ya�PSN��^���߸c��D̎n�Ð�9{#m6����El�)� �ؔ8�O�������7;�V��}�r��{�˦0O�����U5��d\s5f���O4���}�m6Ip���2�Մ�'Z(OL��J!*3ej�������z����f��$èFL�_!X��4��aOk"����.n^%�,]j��[ �EEML����5�5�	����W��`�m���� �kWy�-��@�)�j����:]ٰ��e�2�v[7��t� R=ohjS�=�g7�^1g��F����h�Η�C��́���\9y!5g���q5n�.��7���>`a/5�p�)�A�ћyw~��j��n���7���X� N���ꪚJ�?IzxӺ5>��s�7`u{+�lq���h�d�f(:������4_E�j�zt�is����v��Js�9��	�I۶h@�
��ћ�L(�E�+�r���ڎ��B�}9���9�6��h*H�y#���+C>��=,B�7��i�������~���__g
�'ZDw)�9�����V���/����9ΪF�F�ΰc.��TUF�ݰ��"�OG\���aѱyD��EQ!G�8?�!M%�/��s��,��A��]���V��I��m>۩�d�K{���Ɵ1�D\wރ�Y=��J���Id������6�j@\-)�ϝ�F�/�u���W��ي�+9G�8�V��X�W��qOL�D���26�����ku�Ʒ�S�1��^���&,�tH���j�yXv�|��R����U�����k/~p�xP�!7s̷��hˇ�9������Gt##�����BT����$¬(QT�U�T���L&�7yh���!ce��LH;��P�y$_��D���2��{�|?�m��=������ߚ��;����[3����Zs��L������ D����#��0Q��t�y}�\�2��^^m�}On����b���C���Nأc�h�8J���I�c��`�|�b��>��X��~0���G���働��T��j+|}��ѥ4}�T׏����t�v�uߡ~7��_?9�$ڮm~��H�7�ptU�����M/��w�x/�e�P�בX�vSyy��ɇ�<dk�E�kei+���һ�z��ߚ��PU��+�8*��A�9@�V�^���GT��r�D�v [�Rl}m�@��z<u$0�㶟}��ǚ��|0Ci�6��*�Y&�O�)a��A@��
��6qX>���(ℋ��0&N�X�foO��(�9�y�[2����'�ڀ�ةtn�k�Aؖ��D(�������U��3���Cb|q@���Z�[FaB�VX.H�����gC�]"��$�:_A��h��󟪕1�eٿ}6ȭ��늘��9��Z6Y�p���мy�kW ֿ���g��A��5g���6���x���Hh���|6ǥP[��&^���"H�jK=����3��$����dEH�O@�u]��'�ۂ-� ��|��3�It+
y��+#7�F��7��n顂�91�q�SB���ؿ~M��ߕA�qGx�%��&Ee��L��Éi������bgFJ>�2
�T�Քq��L��AR)��l���$��EV�r�oa���8gNt6^Dm�B�+lL���@��≶=�9f7Z5Z)��%����$�~����c��m�� �aҜ-��+c�m�fk��_6%$���C6��y�˾{"��[<�w:�*��,�k�8ë�&���ʗ��3�\\� �0P��YB)6Q�F�H��0�� ؞�d^��>�jF���o{mO��l�?E/N	����	��M@�kg��g�:������F�S$A�i�;�����ry�MqJM���k�-��)�zG�M�cw@�p]�?;.��Z���M�V�I�$�U��s'cV����z��}��LhV���v�C?ϼ4���L���V2�ЕdqX�8��~Y���"c�)����\��6+%��vy��G:�U���y���"Р�G���T���3/�˹���\�K�9m�D���!�D�N\��-G�'�Y��~Δh)��K�XS������{���x������B��)�P���V��Wߓ���ϖ��#q��LA���5%����܁7 �6�ʿ����[�[:B�|.�`�;��I}˳��&�A�T�ג,�2%Y�d�k6Dd�a�Z":�� X��1ݒ�s�o�����_�y��c�d�Q���2w��
��^�s3 I�I������!��mv��L�q��Z�`��ƳŢ?�zԋ�����!�mp�:΍,Qi낁KtS�����H��#���'�mP���G%G��ñu/������ߨܪł�T��9W�`��/Q�j"#�7w�Ɲ+�%��|�{�j*b6���޾�����GJ��t�:����&�(�`��|a�i֟��������������不�s��d\%�z�[g��΄��x�PXV��/�\`���롬K�����y�(����{�^1a�A��se�a\ư+��LwEi�I%�O�πk�t���D�� 5V�OE��N�u~���	����Q��C���Z.h�v��R�%��6]�z��x��jɷ&�nQm��g��;"g����9:I�+N~q��R^��t���wP�d�ų$dGS�c	�5qͣ��.�u�h�����w�,D����4W�>5㽚xP;o�R��}�ݾ�g�6�������N<(Rn\�SM\{�qKF��<��7��C�� �gR��x��a����,`�-�����Oj���a+��\����l�w�I	יҫ���Z��2B���
V?��_���,�f����n�aq���` �A.���Z��:;,�,��5A�ɶR�����zL��vUbvvm�"u�������L��������ud��gp���-������1��rZ<�8��±��30��K�O���[��a����ڊ�w��W����#��RK4�h��J��8�V���+{rLO�^��,���0����}�%�ʫ�S�����C����fD>�3{�'c�sθi)�8K�Z1�퇯aC� ��m��۱�PH�6߁K?���GN]p�����x!EG����҆Og-�$
�$�T�Ő�$�崣��^O��>�b[�h��\�#��!�t�r�蟎さD�*�^Apkd<����ҳ�"g��N�6ҿ�Z�l��EuT�p�6��*�U�Jx��57j=��_^&�������X����!��0jа�ʐ&���8��&M���/XzdI��В��r�h�#V�&�g凣�8�=��Zj�~�lщ�+Ǡ㱟+z=���2Bл-�8U�26+���f�E�{�/\�]���X�l���0�4~��%^gAj��&Á�l�
��* `j���Vr�y�j	ؾ����%�� �2�������(sg��3$	�+F��:�R���F*�:��
�|Q%mjB�bY�6��G�r������>�=z.
�Y�/3�9|0�qk,P�+.N�.����n���>���k�m���5QQ��ܷ=W6���[���E-�+�]T~���zq%��g�v+N��Q�bǶŎ	�D �����'���(В�;�{羔~��"K�#!����~��Z�[���
�@S���hA9�&ϐ `[���8"�W�K�a�B�p�E���O"(>]m*�h�m1���J=��$��C�u�����d.��F�j�]��_�� ������] 3�#[�e)��%�Kᾨkr�^q,��zϳՠd����ષ��C�0u��?:|e&k)F�&�f�.J:�9_�|rH�����{Z�E��!�e�u�n���� �@(��4�ȨO�T�׃���ɉQ�Uj�,�A|g'-˿�*���ɏ�6�s��-��h��v�c2y-�ٝ������BT����={\貕����/��R|��~U�7|˅��v]kl�4��7���0���U�e�z(?]�ToW��5ם%��b�@�q�g	�H[~�ߊ"�۱�fk�cu"��T�l+:�X^���d��2����j�@o�x���r��F늠�-�܇H�q<�~A�cp��~p֚Bʮm��4Ǉ)\��wc�Мq�������S(�AW�!��$ce��1����?����}�+���������?�����G��9�R��{̙o%c[��P�`�;s5I��Ul1@�e���g������NY�_x�*�����I٠[6[����x��|���$�}C@��k{fUzV~��Cq-��L�p#�|U��X2����$��%��A̍sn3cD⮂�UP��� ����j5U0b�pO�yj���fɻ`������!�8���$�u��H?���+�-X�J�D��3	9E�-��G�.���r�b��.BT�$eJ�v\B��'��G2Vb����%!S�X��ӽ�\�".���|���r�	���AC��֤��#�
�3t�����	(���HS������/��%PO��e�O�^�i�	w;��s�q��Nx�ګu��R|٪�<`eC\l��̽4������&u���JyS̼/�e!_�$�0!Sc�M�M����&b8��;�������D&r(^��C��|0���[x��ZG]��i�q}6Ö���ݢT�%�J*A|�Q%Lp-*�,-�4����^|B��DDCB%3-�ev+M����ή�N�أl�X̗�J��V��f�[����W��b��-�\aDyz��ɿ"�����p��Nkd�p���ai�wv2�8^ *Sǻ����yߋh���:�@�̥��.��� P;���/�@��i�[t�G6�c��s��FE�w���V����A#�x�C�HEm�C�'4�>r�mX{�)P�LG�[s�����֚0:8&j����~ö7]�/��>gUX화B�٨�|���jSn䳎��5%L,<�3$n8�E�m����a}��شS����I���;��<cЯ,L����T�.`���3�߱�Fa�)W��������gu���LN"����[We)���V��=�����R]4�L��|R*Ԗ�$N�-�r�|6�HHD-����:����H��51�J)17�� 0��X�wva��\��K�~��lBE����!L�̊�G6�}�t)T�rA�������7�y\Hۚ^�Qf��0^=��>jz)��L�ž5�v.���a���6�qW8�ԢEhC�x��u�(�|��L���\���<�篧�{}�(�B��Nɜ�ޓ!-�,���4�fm\}lp��ĵW�_�&�K��?�定���5= ah�X�eH@Hz)vs��rT��F�Bf)�xG��I�pAk�N20�v���[�>a�Ơ�d��_��Wj�6B��ǘ�u�'s�ZTԴC�1�'\U�ð]d����p�"��z	�O�T�O�Я���H��3�?DlsD�٦E��#?B��;A�m��i��C�P7�0B�����Fd��T��+v۲�(,N�T"O��һJp��Y��k�ٰ���u������2(�}E�s��;�n���X\�:\֠7�m%ꢈ��@2��]dI(w�6�v��+�L��Zn�:����Pg���䑧��$�-WD�� ���ǯ6f�v�>�E� ��0����I�i�E�xf^����҉�Lg�����	���)��A(lߌ�˦���W+�0[ʧ����%��KP�q�l!�Vi9n�Ap_$J�*�Rv��1��A��Yjh�D��6Z�Z�o\r�aP�wte�w�L����$��0��i`�=�.<�?r�����Q�5m������-jI���@i1!n+{k�h�48�{ �[,YF�v��ǟ�	��z��;������ت�5d��8%B�3&�U�z\���ȑxh��4u�@_ӻa5�J,��9�����L����Y������l�!�2Uڦ9Dr�q�"kt�;�-����2�F�h:<�i�%}�PG4���+�0vX�+'&'�]W`��(�0{�~+���Zm:���"����<|!3���@I�������
���	s�����((�mq�cl
؂���15�Զ�^?-󨣩"L�ep��[�E3��T\���0$1��ߣi/���{���17d�9T�x��[y<GE�`P�sO� ��|Fv��^���c9��O�)==��[%CѾ�i~{=el��u�!����
T�ჯ�8���T��焽	�߶0~ߒ�^�qƱcA�hrf�6���+K�L�\V1\�T��m^�M����Zie��L�**�l�t��k�g�#j9k)Zx3���2��e0+��Z�m���%h'�(AT�J�j7/�g)�X���J�ڹ�8��٥��.e*9W^^�0K^1w����I��n�a��PS�}�f�Q+@x��y��A�����D@ ����D���fi�:X�$��$E��b��x�0�l��ȳ�&���P��`��v@�h�>�RU��� Ӿo	C�k��ӲG��}Z>P������eYbt�6I��Vm��\��T`�fJ��B˺�V����k{B{*����"�;[Xƅ��@�ۭ:U� K�܃4�J��/�uK�6<Z�.�Z{�{��g���U�<���,��4�u]y�H��6[�f�|��*f���,Y4A������[�H`H�'�ߥ��@��aDD-��r�K|Iv�*KE���-Μ�<Ri�}��q]İH�J`p�%i��R�5	?G�g<�/����f���j,� a�5v�kYg�un�j��"�v�t��n(�[�E8)��%��K���0!-��Q-	@�/�YuQ�d���I�RM��(�-�"��S�K�|��=>o�2v��2��kE�=�s��_�%�U�"�t�L�(mzE�����g�!�Y�H0�z�ۼC����I�"݌�]�1$t�PNʚ~n+/�vUшK/H0r������/�p�9_��H �̪�sE�|��+T�g�Gu3��{AS:3�%6�O�=0�\0��t�,��C�>��V�&ܒ!�% H�n���������:�s�ߐ���Ri��Z@e��4ݎM%up�,Ҷb��p�g��jˬnj�>U�}HiKo�ӷ�ퟱP �O���;�:��
�Ni�BbӘ�;?�{�
H���c'����ux�A�� �3��n�{�!"�r�`�Rh}�?:�g����^7j����Ku�YELgsw��-N���[�{���5CKX &I̸t�dhp��C�XpH�k���4�O���<9���D��,�g1��K5�;�%1�7Z���\(i}�W���rE���Q��v����_��o>����|�x=1��l��)�Ꝁ� �Ĭ��u��y��:�#�f2ER{�X�T�ۆM)����]R)�HJ�N��W�;oy�bD���pmE�9~!0i�ޘ����8Nx�l�*v6�l,�WF��zg�FTMᯥu���Y�0|�{U�	�:�$��5Ҏ-�*��O-��X����x�qIP`8�d<6o_���z��ƠO�
��
Z�����h��b�/��Ӣ�O|��s����7h��  �1�P�7i��AY*FP	�l����L���qF]���w��6�Hh�������!�S?'�&=p�!��rMPV��q�+�߷�i$�v�����N�'���9�騼�;ԃ�Ͼ+X��2���	){`���1�&rw������<Q믋�ᨷ�Bh�|��ΪJp�L�?^�*����Sl��ju�<v�W	%� C�h���I���$Ɗ��a�Ь9��H�ݤ ��tK�}�\Q��E�#]+p5�31T�� �?k!�`�l�⃥ 3'J�&-� �$���`u��
����P�n���IPu���)�$ƣJV
-Vb�EO���M���n'|�O-n���d�QY�d��EI�5*�d7�iH	8��7��E=}���&J��x�I�O�zF�b���*�������8�a��"j����uH/��`�oN*��UN�0�C-�x}t��Ԗ���w��I�`����:*b�������	��v�G��˾5Ӭ^�D?}�9��K���h��=�rN_������$V�����`~az]1^]1E��Jn�a�i�u^<r���s7���#��,J�����ĝ+��l�T�5�ꂦT8T~�_y[hkv6�-��7�9����?���ь"-�g�i@�ą+1ؾ��G����p�DJi�1 ����q���
Z�5�d�1�|�=
���[b��ε�bN�]���7G4u(�ss��{
�xAc��sJ.��}>~�(��56�̇�3Y��Z7]+�7���ח�G���@t�e&���c2�K��MŜ�좱�p��Yl�O�ڱL�������r��pKj#��T�_2�*�1R(���O(S?�E�.��C �,���[��֠ ��wMr�Tz��:r�M,\�9Q�q�
�\n^φ��;3@�l�d�W�
�f!X����(S�C�,�lK]��[�X��D٤���n�b����W�;Ϊ"|q�?q�G#FΚ�e�e�a(��d�?�汥N�X寧�qR���㷱�����IW�����t�5�ܤ�'
��0}�lDQߕ$K�M#t�gD�.��~;1��b[T��o�v��k��_�Z=��ߓc]���ñ��������Z��>:b�-F�\�^��;jm"�;L�N~�F�.)��ӈ}`��([/�JN" ����]���uM7���ۚż�h��R�w�a@t���,㶪��x]�JA���jn3���ԛ��f]TqF$���=�]�JAޟ9��椬����F�~�}�'��\A�n;����ƽE~j���?ֻe�f���n(��U�8�uq#g鵻Д��
��԰�H�iS<��D��o����.ke_h����GQ�ЮN��0�5���n,uF,�T"��RC3Z�/s	Q�ƛ���4����F�_��Al�R�+�Q�ս�u��[��o��h+T��ȞK�=ҳ���)�f`51l�W��l�|��W����yi�Қ�@ȱ��y��/T�e����T��!��0���ǳP�dB��u��'-�2�%�H$��ѿqL[4�[v7ѰnUF��U��S�3�P�m���E_^t�<66�`��0��.��x��91p����VQ�����멥��O�!ˠ�,)�10Pl�<x_�,=�	k�nIZuH
ܮ�EWj�����m�)�Eڅi��4!�u�v2�N�/�ٛʃ��V�4���P3���N�h_f���D�e�ȎÐs	Me�?XwGps���yF�\%��f�\C�3��}�����d����Q,��5�z��2��xt-|��;"�8@FQ�/p���9ɃF~0'a
g��{�BQ��$��-JpM
4�� �ֻ���h�8x:�ި85ݖ�,z�R�آ#A�(���>c��k���9��Vk��J	�OY�mz�Jɦ���P:��Le��A��]@�N��Y����Z�9Q��m�_���0��=��v�e�Bl�{�$O��N�M����B����i�uӥ��`~&��8��f��}c�u��NѕF�+vL��@#NY��/�:�v��/��gcjp�����#��68{��P�ùU���̻�c�w-7�W����0��~��P]�����+��1�f{V.�!�MY�p��~)@

� ��:������>��.�)�Ч�0?j��R�yL5�emm��;�i�k�c	Ϻfq�mPD`J�����\��ʬe�a��Y���8�hI�QH�o�t��bN��1��@�[�.�,G�,ݚ�d�����]6D���|JfR?CFGu�-qAx��i;�����h	ĩ 9�l"�!n��'�=C�>�.%�E�|�c3/Z�������]�'��+e��>/Z;�"��=�y]��4S8�������ޯ����6�+����b�I�t����ւ5���;@թ�Lϐ�x�`$l���6�x�d�I���wl����Z�G\��^��^��8��=G� ��P�'ݞ�p:�p�:N1-�?	�1\	��B,I�,.��{~!�"o�{������;�����*e.
�+�)�UA'X�n'����<��#IK��0����a��6k(�㧃j�go���`��7�ۧ��{v@�`���ϓ�j�ZQY��5��Mbw�fCL��":;$J�l��N�yn~�Z�?#�25�6�=�8,]�6lP#ݧ�ڹg0��HZ/���0.�[\/k^��(PR�J)-#̃D���3,������f����`�܊PUI,��?	�;N��&Im42Rv����Yd���)FՃ3���V7�FF!�%UU��>�vOL���Q�g�M�2��C����J����C| k�y���A���� "�����MHB=���\�#�䦾�(:��MfW�u��g6Nvb�L���[�z�ޏe����_���豼�8���dދ;�u�c���<P���eC�t �L�mz��%������0Q���!OS
�~ÌR�ĕj�4Y�s�����ŋPx[d= )��,�]����F�024��0
��Ϛ0��]dǂ�6�5���5LU��\0��Qo�B;�+'#}J�^�iN2;L��m�A�1wT��J���m32xR_AX�݊�T�>N���#�o��J�E��[�T ���\3���ivto���W��=ܸ��=��-+�	���r,m���R��	�������\���O�o����h��fA��?ʧ�,iQ��*j��l"�Vgf ���LH�7��U�9��o�yKb�E9-�_v!�st�Rٕ��}pǼu�J�F�$���8��cЈ�0�q�L�.?�y���9T��	D�u�x�b�¬�o��`�Cv�_�)|�E>g�a��������ݜ�aKo�Ƞ�:|��G]j�cX o-�<��Ξ�'aK�o pM��Q9*��VO��S�y܄�ց�
���K,���N[a'��ni���Q�y��\�b������H����~@��m�%I(�/a�88��o��'��^�7&�vzR'È���G$�e` �Kw{�S���?��2��O��5K�᡾���Ҿ���F�ꛑR�W��<��;>˳����x,�9����p|���W�w@��(���x�-�'L{�+�6+J�����8��Ϫ���eJ�\�w���M��d�U�;��m�6��J�]��Z#�z(�Z�y��Y��+�H�¶n�r�~ <xDO�_�.U�i���Y��ܝ��Wnmag���v)���)Nt�U �����l+��S�����=8�S��,�
���s-�A��E��#=!�bm�o��]��#������\�7'?���tO#�jV�#V ��xq�O}�d<z���	8IF���`�]jrkL9�n�Lm�@�����.�,�,��H�-VW�C6�o3��V��cG�W�m��)���چec/�n�G�Ο*)����^r�ҭd��8�>��|PE��>;��"�X�Б.cȸ7�2�&�1��Q!���/�ny��P��|�t$�̨|��6��`8\E0ݝ,��,��d�[�8�:��X���SB���Q�&H9O��o�M�DMP$u�eF��k�@#�?+���M˾E�c�/���Q�nceC�t��6��h�9q�|��@r"�3#���X�\�=��	���۩L6�%��V$�2nӶ�a2�Q%�A��y���F2�#��)P����t�{��f��	��� ���MJ`�7\\��3q��Vr.�f�G&����JR�W%�>T��5M��>4�Ұ��g8!q߃��}���G�[$X/m�2�.#0�;j����E��?�L8�P�	(][�2���X3.V;AN�3z�<B�Z���\R�EM��,}Uɻ����I~�af��*���]!�Ғ�,	�U�X�Sk4�jq8�}���:�i�d�T$��]��@��4��Y��[�\m�0u���C�h&!��X$]i�ȣv����&�=���O�7%� u��{C�:���s~+��ɬt�i��Q%͇{�Z���kfg;�s,q�v<E|oz����Ʈ	8��½rW*�}���f�=���)-��GdA����f3t�y��i�]���~bߓ���S"D�	^.'�ݠ�3Z�K�e�:I6�NF�*Ax��(��/&�O;�H���%5z^�۴'�n�,-�1 �]`=����ǚ�o���B�D*�tKF5az����v����(���5L��2���XfW���u�tN���>��*�ۜ!�3T,�K��#�3Jp"s���H?������P�M������*�B�]Q4(�n��]Ө)���n�Nf�W������M��к_�
��f���:]S'������ @ ����/�Q��,lj2@�)9���a��q4QE,�u�����f��F�Q��2�bj��Qܠb:�宀��r��q�k������rmg��[2�l�-�3�cڷ�V����@���}���a՗��Z������~r9<�9~(7���m� �~�6�����J]�ѩV5F����]�V.ժo(�g+��kp��*�㊹m/"y��?5�u�n'^1A�TPaF&���0��Z����]�6��h���`)p�B����_|lA��"�ф�c|ּt�f���g8��Ӱ��@���!�	5̳����|�R��z^�a���ս͝l��)�������z���:����t��$�!h��}[�������֕s�m�#I�Hy�P)�p��&TQ~��4���6�1�c�CI�+�o�f"驰Ԩ�d�~��xo���9=Km7��hs�@�@RL�_YU"QB��Q��Ő3A����i>��������!Z���)�80�v�B�)\B6p��S��3ё�^x��Q��xKx���M��ꃃ�*���_�����iD��Sl]n�pC�3-������$@��qZ�����82��/�<�h1ڪ=������C��5t2���N�뽕�+��/�f�\3�F��|U���}M">�ί���g�L2p{��Z�����-�LV��L~J�^�h�i0^8� k��AF�6�N�� �,S�ZΊN�H��YE�Ji�b��0̝��2 �P�	���L��3��eY�����&ְ5q	h5�ԯax|ğY���Y7�[� e�Z��p�R�e;�%�R�A���z��^Ց���cs�Y�{��?I�:�[0}����ٌa}�w�\�.1`�F�SM�p��l��+�5*�Υ����Z��������Wf ']�w��-� �����;��a& r"�t�$�r��g��1A��9���Z*˵c��g��ʅdL`��P�f�	��_S��^�5�g��9��H�h&U&�x7�,��[����@Wp�\h��o��zS�4j���ͺ�T���l\��?�bq�5k8�t32iV O�v��÷g3���F;�Fs�����{���I�x����~�����}M�_�Ђ�����؁r�#�6�e;Տ����ac(��$NtS���6�R��������c'������h�DH�d�BRf�tAaޫ�r�F�ug���M�M$;�����v��L�r�-�)����)�=zwyɟ���n�:F�#��Y�	ӻW��et�EPNSI�x�F� ������q�w���GS���t�٢�nt{7���b�����3����Z�A�1e�1 x����t���@n޼x�k@b�T���� ���Ho�UizJZ:%_U}
�0'��MRS(29�8�OiRKɬ7_�p��h@D�����`:��}c��5|�Ot��X-��!ķ�D]��� �iъ��
��oIy�k� =�ٻq�?��@�X�*�� �Yd:���=����P�kRpRx]N���j�*;c�P$����d��Dؽ��?�T��3�ZC8Ư�����d}���m�C��}Lew��z�T�˫�W�m-?~|�)�ߞ�
�]]0�pH�I��-��"������q�4!LiЁЪL>'���ٯQө���)�J�u�b�m}��7d��N�s��_[��75���W:�1d!�������x�/O���F��mM�ˆ���1\��Q��d@���Z�<T4+��;�~��)/TL׌t��<��):4Hm�H`����SG������|�PF��d."^��VW֚���(�.^rP�`S�,��Z����Z���Qր�ƌ�=�BA�*��M�*+/��T��sR�V�uB��S�o?��$N/��RD`˄����:]X���m2b���J\R�Y�p�M�:�ȁ��⬭�F�{ h,���?����rsf�_vA�(�k�A�H�5�wwvg��*�g"���,I�~� A��������ˊX�Ds্~h���l���7f�M��.!�	ca�ɃB�S�xP���i�̦��]K��捹gD�6��.�8�k��
F�UĆ�j�x�7kf�h�t���-�p@�zġ��] ҏ֣S왱e�@m&FT��v�W�Ɉd�rͩC~���'qr�Cj�S����a�0���Ҋw�C�ߤ#?�$B��B50��婍z8���~m�>ᚾ �-0�UEh�	q�f���z�kiɭ(0NQ�zO��-��}U-�w*H���H����M� u'!�/ɇ@��щ���2hUS�G!j�L>��J��s|�Jg?(j������� cn�:�� O���	 ���Z��	]p���t�z��{��K1���˩�L���xd1'����*'.{��E�M�H���B�����&ן��A0��"����W�/=�\���J!N��&`Uc�W��Ya�X���ir�wȏ���7�.5~ˁ.}���y �f��$���|�<�{YI�\���0�S�W��{�s�8F��h�7�����N.rǮ�ӕ��F�d�G3����:ݞ��a�(1��,j��į�<rz4WDwb�*����M���J|v��4���=��B�6�M�en�?O�vw��3"%r�\�G��6��\m�b�5����0�bt��L�)��An��)�	}*��l&�w��!�Te�BJ�:�hǒ�u.=,�и V;�B/g��f�ү:��sh$%ۜ�+�I���gu"�a�H�@��TzH���
V�bm�RM����{�xη�E~�.�0V�M` Q|[���읓G)�(���_ ��y�.o�c�fȝ���*Kʅ �W��N�������(�W �#Q�tr�G���'��s����^�j��T���Mnɱ	N���B����$�FÐ�G��`��0V�L�e��D`�V�����5��d�Aԅ�����V�K���Q�#�6kt#"[ ���nŠɨB��K����l=�<{��OU�U�^d��6��#�r�81܀�6�!
{[&s�g=�S][��^�iy�� ]�V���ka�P��z{Νvk�Z��1�-_�t!�i\C#�W��P�gFԕؕ�Z�$��[���<8�v�g�Q��	��c�n�����{5��zH����!f�"'S/��u�P|�ȇP��J�Eg�������C~��ƤǬ�2˞���*�`h��y�;�I������ĵ���7��s���x���`%s��dFq�5��2C�H*ZQ��%��^!�yHɷ��/��̙Li��F�?�آj耐k�C/]7���Q���&6Lա`H�k^ȯUT>�D2���*Ʌ�٢W����F�ˮ��v3���,t��#f��0?Z5dy:lB}��X�a-�+y"М&�p�������U�o���7��6��+�8��������˶��n�5��_�JQ&1�`#�F5:��]��qy%��5M.b-�=z`YE�?sF�:!�8ҡ�zq����a�&c��O������(���f�]^@w@>�$D���j�^@��5e�8p��к�+���Ǚro�M��_rtͿ�w�����{�A��c�o籥.�@�{7�Z)�h�Xx������8�Q3����ˡ
�"��7��:ۑԖ0`�|[��} |J�6���"�ɷǳ 5*.X�/�y}׀W!ɫ�ʔn��Ǆ�)�t��c�<�E
L��g��D7S��?�WҢz�)�^f�V!t��CQx"v�e���w`���Z	�aQ��z�Dl������.�����)ѧ�?�.��wy��z��^ve(�%��O5&XD1�88@ -���m �pZ��c�W�N�Ӕ��JD��)Q?�N�9��'03X��IA�^ڠa� �⁞��2����X�X𩩘�(r�l�]]����i�C�����>�j��w2
�LP��kc�m5���R5�V�sy�s��D�OX_�NY4��ur �&�lAo��k�Y��G�@.SűV�x�b���/��mD�y� Ʈ���8���3�y�P�h����c��E/����-d+Ba�{�@�	�/��?�̘
x@B����4=�D����U��{��fƦ�k�Dl�y۽�/�J��䇵G�!�CY,7�m�V�St������M����4>↜$?�[��ƃi����IrN�§�6�ʊ���c�z�W=�"r��(��l��\Kp[q0Fi��U��G��C�6�'㡝r�H7GN��ZgE�k�E�_�V�͵ĪsM*����M2��{&$~, ��C���������ЬG�>�|V�l�ю�}f�oֵ�"��۝��`���R��S���㽭�*&�@�8�t1(���;,�J w�Jv�؉d��iTk?�]�Z 3���L�
�ʓ���=�!Kה=$
j� X��:�th���Џ�D�S�����UM�"�0�W��y�͆�A0��e��x�
4���)G��=M�c��!{�����ǐ9z����:_�D4=&�5.��m���w��I�i#���ZΌ�>��iԳ�"����m��W0 ���t��۰{냁#m�M�n�`?�o�����Կ��U�e�`�:z��5���� ����.�	�S-�)/��0A�P(�UC{�n�Y��{���xT�^��O�Q�[�0LwY�����p!iۯ����T����������a��=��|�x����-�N���3@�x���cM�RöY=��U�7��joQD|e�L[��&K ���mS��(���+���}�"������<ae�ݱ���C�Lz7nL��7~S,�V:�� �VnmC�3��b����_��ć(��eɋ6E�*i�/��W��MܺPj8]�Q%N�g��U�<�-~�2�����/���O��	��THPx�\}Dj[�􋉑�ԥګ�ߠ���[-��s�.�:�)��*�qԍ�>�*[;�l5%�<1��R��~�8�
�v�uQ��f�x`�E5�Ⱥ��H+����pe���*��c[�-�A[��5�+(*��ʸ��B�K�^�/�(���S�i}�đ�"��ʝ1���}� �:�-�.ߘ$y�H\䉆�;�v�^�mjɧ�NÂ��[�|���8(�	��CF�Hٲ��n�8Dq?���¨��p4�m�:��7<�
!}w#�g�?Z�O��$0Rem�C_;2p�-n�MZ�%���HWE�}���Ͳ�N��i��H�U�6\�"^�P�.�z.S��Y��E�ک=r�"�؇b6^ٙ|��	+�ǘ��H�mE�6.� ��*��*�Ω�lw!:<���
>kO%ZF�cm� ��V؁/���C���N�6@9P��*�Y�``L.%a*�=nL�Z"xf��� �~���|~�>��_�#�Ush.��ł�	K+�>!�9��a�N��zB�"���:���ͯ�u쫯_Ar@�e�
�e��Soc0���<�rhbu�U@�!lg�3��3���GF�m�.��[�u��j8�Mk����ܧ��vc�����4U�|����N|���t�t� �i*�	3M0�<�y�EE/ ��>��F��{+�| �݆�}�z���-�FX�B�`�zϞV2_�1q�G�-�gn��	��Ԭ��b=��� �UX&ƪzlˬ��]��K!�;.��B��z�'=�/��W��E/�He��iu23�p��aa>�5�h�X2g��j��#�R�{���!����9��Y��Y_z'ȴ�m�ؚ.�n<�� ���:Q���n/z�i#�-E��iZ�	%�/0O���i����6'��K2�=	O�<]SR]��nC��~��,YYQ��<�f��SoBﯴ���G`������/���G��D���7eZ�V<6�PtG�:*��1�K#�W�?
�H�[
e"zI7R����1�V��?`�W�@ N4�i Y�r\����Ĉ��U�}g�+��p2�E���:��f��q�\�_Ɖ�ЋG6�E԰��ٱ��P����w�.U� ]T�_���(�Fdi�����/��cL+�����B�j@�l+_Orfr/���'�#��cp_��\�<m�A�RD�sm��S!U�nUE���ț��g�c���F��mp\��t����-�.<��\�^�4��g��^�Ozh ��E[v��Z�9��{K�����]�j��;�Vk:ǁ���g[��G��5p�̑φ
�1���f��=aI�h|Z�go����uL��Q�DS��vi��F�T����ʕ��( ������!���{������g�%�'5fʴ.f���'�#	4���kɓ���ۋRiҕ�e���X�x����e�G�?Y?�� }���^Vp�!�O�a����X`b���n�2awﷇ����Ӂw�?rEwɄz���=���ɕN�UJ��ܨ�"#��C�?�D��;����bɈ^�^�2��dX,�� ��Ä]�
�Σ�phQ1ͱI�q	���d�4���٫����w#�F���z�~䀜���`��S '�`��A�dbJx�ו�oX��G7H��T��榽A%n�d��3�E��x+������݈g.�V趽=H��x��:{̮�|J1��� ���C.�LȊ��i?���n}-.�KJ��8�g�2��n�7�d��8�� ?�V�K���p�49s��~7�=� ޗ]�.��ѝ��K���	���>�t_�M�3BvZ����V)Ȟ�h[)`�	m�iMG8�7Y�E�l�Jѱn��]Tw`��,�/ �\��專f�a�]��ͽcx���.ţ$G�|Q�1�1�h�J	Tj����T:���[��0�|�h4r�\H}�댖^,�t���#�uF>��C��b���S���Ǥ�Խ+c�����hL�;	��z�2@BL��n#�̀s4�&���_�;�8�Hd�;�����m�����`�"U�4���r/ef_�z���O_�~�����=��]#��3(��u;�hQ��2��1�(pUb)������Yjz�Ӗ�� Y��i|e*����I�z��:�m�c�k^�63!�,TK*ܽG�L�2�+�n�"T���J���wN}I��ɐ�6s ��sN��^ ��X>�gw@��ˏv��h�0�~շE�'����Ձ�M^3�䅲�w�����HwE�(,l��c�b��=ؽ���[�:A�Ig���Ll���΋Օ\9~�w�'K�P��ۻ`!�'��*x�l��X�����"�D3�4	UG]1��S��
����&o���'������q/��Q1=����J��z��y�PN��L͒f��S�_����:��;	��^=�����ľ���@�TP�z�&��������Jbӊ�A"c��{,$���Ѹe\ �(���͢ ������eȵ㕂+?Thv� "Ť1s��G�AJ���2���}�x�����c!�:^l+��k�*M��1GΓ�!���+�v/\��FW��E, Ԗ���ڍ���{L��4��V��1����:4����ys�1�
J=��}d��~��Hg�+՞ҷN�3j��i��`�1ź��K�<�`����Z�3�'X"����Ϩ��[�ڿ��z|:��
�����U����E��x���bD����jl��%;,q4�E��~"�h��t�Ɏl�}�qs��Ç����[oo�E��CV�����"ܗ�N��:L� �x���E�a9�l'F.3�;��1���rY����Y�n�����76���#X�(7��d���x{j��:3�#.�.X��4cZ|C���0�O��ؘ	7�*H`�&�#�H�.<{\��o}2�t�T��)�.rLIű�����'�kx���\�.�ˍ�3�pܽת���4/8X"po����ؑ�1�5��\�U'܏%�L�}�Fˋ�F�������T˱�x���$-�����k�_��$����N�G���qB\Jr�%��R�Z�ru�C�BӚ�%?���W-=	gIlT_�H|�����Q��H�.��bCUm�GK�O�;�2��v�:��y	=�l��لo��H#=G�h5���#�8���#d-Z��mrH
D��T�B0�Dۂf���yTd^F8�E�,���.�)�YX�� �w�7��sCƗ閕�\�K�2p%Ix��.�U�Ӧ��Dn����u��ܒ�w	�7�CH����zs��l��pP�Tm����a�����!!��k�:A��s�����E#��c42��r�R�S0H:�xH����o䀇I.J�4H���8��P^`2����v~�[Z��\}aVxn%o�c�r=��5��E���I'zm��4���m�{ ~69�Ř���/Q$���'�7���J�#~�0���wN�	�9!D��[;��@�J��U	 d ���*f�#s5ƹ[���~q1�v,'��>�v�OB@%���{��j��Ya~�ր�ih��ߺI��r�ꎧ��O^�и��e9�Z&"��*��P���e|3S\8*���t�z�M�j�j��D �vƉ�����l'U�N���v�=Q��I�ט�m�x����W�0t˟�Ϳ<�a�lV�n/��D.��Z��VY�f�Y���8��P5.����s6'&�<��ƺ�z1�`�#��ET']�7ӹ(p�D���Y�輤_p��8V��c�(�;�9�Ie���G�=x#����ѐC3�G�UY����LJ��*��C�-сd{��o�
��mH�b��g�ѺM��Kμ��9_�2������],^bko�+9��2�1��ӧMߨc��~TK�]��9�� �<�	�b_9�ER��~)�Y��Hr�_&'nx��/�w��C��0�b�RnZ1厧w>E��d�`�@T���n�@R���"c�J$�քq �(��θ�Y�Ekw�V����LLm��&�z�,6��j��b�~���D�1��;�H��*'b����g�r��r2г���9ǵ�H����XQt�8�)�D5���ҵOX���G��k^s��|�k��d��"�� W��th/�J�R�Lل
)P��Q"M-ƹ׷U�����+�e9|�/�A�ȫ�2#���ع��$�>ҷ�D��G����X�QF��2*�fp9=i��6ӎ�;&����:�?�fJU���ٌnyi�,�N���(���m���4AE֝�Z�~����f���O�"���2��j��z$�!��eD��/�]�o��Euwmn��R�?�-��uu�ݚ�87u(q(_*R&n+ X�l��o [8ۏ�-柋a�����s��2G�r�v�>0�J]��UGp�c�x:mH�e����0&���X�3�����Ғ��e�WҢ��ejأ����H��T�1��k��D�Tf�V�Fj�wHi�(Ay�0<�{�H�`���LC��	��u� D��i��$�?��A��}4��دE�[Y��L�CC�$���I���0�rۊk�����}~�9�ݬ^}+Ǩ���l��2�7&�$:0Y'��@�U g�-��{L���u0���J%��-�6S��hߐPH�Z1��kIHz?}�i��PHc�g����m(t6��Q��h�r(o�ªf��4�˒�4"4�����5�N|s%���+JzAw>:<^�K�Rd9����"(T���
E�b���Eq%,��ܺ�=�8`�eۃ�2���+aA겤5Wؠp��?�<�F����8�$��=ضM������/HAm���ū�r�%���IS�%�ُA#^s�K|�U4~�>�+N��B��sF�,7bz+9��ƥe�&�	���4��h�R���
&���C�t�u,����Xe�����^��gC��W�yF|��bDECr5� �[i��u��zn�������p�CG�~͉�P0���m�o��3z���h(z�ӽ���_l�範t��$��)�ܒ��$G�:�7���7h��)����΢�9���;�ݎW��Q�>�`r4�Aaj�OZD��@|4�#=�EU�������d�J0�$�p�a� ��<j��G�4E��r�w�A �/;'V��Dq[��X�B/r�t���x�ݷ�.o���-ES�U��Ǝ=|�gm�t��l��Eb��[�]L�\��q;�=���2�A�4����	^��$!��Diˠ�/�!�:�)G�l8�ϕO��33[��5S�P�I��)���|�@3B/yq��4��Yu�Q�XN]�5s�����m�UK�B�e��6�3�P�:�Y�
p{t~��z����2PK����+�Y>`i�2e�\flK,�a���8N�h(��KE��G�B�>��	^b�Z*�4�Rc'�}��2��hߡ���:pTs�B>zʹ��zjO���2�	��2cB��͠�j���ojc�u ���O[��j��E ��}e��8a.�-5fI�ʰ.� ��KŠ�6�c�;|���X�^_����Q{�m�	�g��,�l&�H���p?zN��9cЦW�<mM�~���Cc��.l�E5{2����M�A�'4��9T3;fX�BT-C(����E�VBM~���<�	�aX�����>�jD'�AvS�6�p�lښ��琧�a��o~�Y���.�=���� @nF��f��xwL}S U@&���R�����#��O F ���J��ӿ�Drދ�,D;�쑿nx��&��C�TwE2��<����l���scd=e�>�'��+�P�,��H���5=	�T[#~�&��5T�]S������" O�T���ހ��B��PaV����u�.����Q[[|��fwZ ���aiZ��/t�I��yrWOaW��c�z�]J5�T>�� iLߍ���-�y�hqr�������#;�R� #���!�%�t��B<�+ &���@[$�uՒ_�ƻ����
�D�2����E��~�<7B����`�Z)}L����;kӣ�'aH���
?��X��LZ�{�_P|n0�{�8�����bLy��Y#AX�@Վ�M�Q�3���]\�bo6����fV�ML�R�f�m<������Pr�M���ڨVLb�@������np�Z�.�Rݏm^\ů�\Ө�A���]�o?�;��Zl�n��|[$s��x��I�fJsm�ƹ��+��e�5��g���b�Hԛ.�_	;�POQ���F/� ^K����*XxfKP��Hw��������D�+Ԓ�i�o��m�ǁ��T�ѣ,�A��*�� �������;,�ӭ���!Kv{e̔�
$�IT	� .�Xi7��VZ6Y,6��i�n�.��M6O,�0�Ӓ����=��z�~���7����g?g ��U�a��D���Ij@���`����;Ѧ�Q��aߔ��Q-�&���Q	�H������+)��D��.�i�=B�5��Y���b,��lk�+����W�?o]D�%����x�&oS{��Mֹ��\ж�ꘐ��"���=�����w��f���]{m(�����q/u 9��]�vlv˂��bd���`�n<*"w�6�RS���i�Gi![y8vރU�����J�1O��y��n�;H�[���	��J撁䯻�����z�$��'���ɝ���s�aaB��b�4?���6�<o�o�3��-��w�~�2�K�Os(z)-8.4���k�u�cw��dJyo��E��j���ƔY�:�b�J����L��j�К�o�$A��H:=���2B������4L����\A� |2�fWQYM��b��'��C�/�g":�Y���C��8�,����EX�zlFuo���]E{L�"�'�А/���zx���h��a½}�0$7F}�nX�v;x�������>�#^<�����~��:W�qe�ܞ�:���ˊC�ԕEv���)W��|�A�����$d~��l o�m�Ԓ|Q Hg�y�nYN����Z�R kٻ q��g����Sa.l�:%�PZ#%����* �� �q�	�F�&�.��|��F'��驕�/D��}���\@J�kR*/�L�<���/�#�_
���{!����x6�mm���-pgw����J2����s�z�a%X��g��g+�E:���=�4��)2�z}v�X�*��[&;����:�2��u���T:�W)�T���q�*�;.Cu�x�ۑԛ���%�y�(�ژ�\%���X~�Xy���S��+i�2���Z�`����p��δK�b�:x>\8т�󮑷�s~rihKnpx>���օ���!x����Ŧ�'�o0�xC�0�A�u鴱%��	�����2�K��7�n^@eh֋@ZNY�W����{��n�ɥ�ʌ�bqA#!T�EKk٩v�F��@d�+����&����k��p��S�u�Z�M���I�o����%��>y1����!aB�����ʹ���	16���\D�h�i0�/��k�:9om�~HC0���T��A��p%I	�#�&��w`��n��o�%r{�zg?�����_�?b!M���Ǒb��A6sВHy�7��K���>e;;ǵ"�a�*���:J|��'���m�`Ԋ@A�}'*K]��0և��������3|���6M$���43�*�	�w�OP&��!�AA*+����Y���ZRL�v[up�x�vyT\��iȠQYT��j��N�3=g"\��%ט��$YƘk�-�8m�}��z-EC��q��/&Ҏ��V���"�ko�?�nou�m^�9�V��m�-;�jI���#^�W.`W�j'�A:Л��z� ݝ)�1V�:�Ǖ��ɃY7ӄZ��tȾ���f�/�T'��rZt�K�������bP�W��X~��Ӂ������E��!��J��;��/��Cv��]�S��Jq�/�6�h)v<Xi�����BF��`ν���H���v��JL�h� I���Xb*ۦL�#�;��B�v�^%g��	6�F��m˖'�]g��om:�$Ak}������):��<z�Ϛ�<AHl�-nF�t��$��R8��w��HӦ(Z_�G�a�V�k�a)B��鈾��T�'���6��q~��v��w�?CA�
�q6*,�_O$�0l�_AY���k�;	�/)�tk*S�Y0���I��T,R�W������)Q�Xu������n��w�޲�Ʌ�hZ�Ⓐ6G+�\V�k���%�<=�8�;� �OYR��Qe�&�)Q��F�4�wW'q�<�$Cv]��S�:�sC�ŏ��cO��`�������[����0a���_�w�ULz��P�!P��
U��3S��B1�o�S»8S��{�j `a��\�-~D�M���;��Yy{Y���W=W%��zL�G��P�I4�v��9����y}YJr���oˍ�[Q����D[��`(�MSǱ��w��r��#�ɉO�Y��\�3sv�'�����C��0�E��,JE���DnW?�����C��e��v�Qʶ.Ƿ~O��(��b�t:�q����L���*����/��:N�f���8��������;5]H�W�N`;u���`�P��e.�e_�'����<üo�}��0d�Gce�*�'��&|b���P����Jr�KC<�%�A�`T����M�z�ׄ=$Ⱦ��?;�Y�4]��]�+&r��$�Ɠ��|c�/���o��=|"@��qT�o�C.�`���я�����R�Y;6�^G+����%2�'U��I&� rg�/�5�8�}����F��'U���띶���5�A塀�Q׽�X���M-����u����Pb�]w��E����@rht���F��9�gr ��9ó��	�s$ ^ �Ѷ�{#��~��T� ~ v#��OmVV�T�A98����`ǯ�~8yE���B���Tm3UK�Ԩ��$B���O��g��6`Cr��B{�:��4E`�a���y85CcguG�f�����>.��ˣ�	qc�쪚
Շ��7?��c����Y����";#H�:���V7�E�����n��q���1�,�N�q�#4�k*$�㦝�����݄�a��@ �k>T�}l�J�W/.�4y!׹	��:��X���A�l���Hs)�.�/n(���*�ǩ��%�I^|���/��L��cxn��U���e���C��Y��(	��<;�x��"z^�W����FU1n �Ȯ�Ӈ��FOv٨q5�vtS��=��tW�h��"X����sf-�ΟW|���l(�1N1��s�ם ;��N�w��1����T!�1��G�^Ǹ7� f�EV�ƾ�mE�`��u���j}�#�gKAYD�Q���>l�<
�}Q���89��y� 5��7�*�ͫE-{�\�^�55%D�T�A��F��è�Ղ�
�+/X�g�t��z�)�i���yY�R�ny!�q=��r����*?�C�5H��+�����gg��]ib��0�
�5����؞��JB*P�5��;�D:�C���F�W�[r�Ee���ڰ}`5���C��L�k�4�!��ވbT {������1�ݤ�|MPl����ٴX(W�t,m����h	m� H��O��T��;[��E���A����ua�7&�b��5�C�tb���K�´�Iw���䮽��jw��E&�gh'OM�:�-Q��2vG�%z�m|�瑨,zjt*�`ݴ~�Z�I������T��-�NR{�HU��]����\�;��Yz+'��#�%�D���/�LA�P��iE���l?L���b��\���UCi1���A�Ђ�T������CZ�[c���*�Zb�n��_�cl���N�(��~X�yT
�ic�~2��<I	�~��g���7��3�a���؛J_���=����+���^�6U�4|Z�f&n��0ߖӨ4,D�@�^R���F�o]]Ĉoq�"7B�o�	�v�Ss�В��bg��
�x։j�/�4���I�� 0
��)"xtޟ��uCh�P:�{hM��@%�U��7�D�n�!��� oG*4/�O���vۗ����?��W���f��^`�T���cؓ�MTX�P2�_���Uz�!�+��B[��#J�s68<�G������6�<�fg���M������Bꁣ~���@��Jq W�����Rhj���.���T��e���[�y���Ǻ �hl|d�}1���t�J��<�'�?������D�<2 �Q�НR ��n��|�ђ����x/��y��YeBOۤxV�ۈkǐ.2�8�N��X�|��{
'��K�׆ ����=?,�С�K�
T����j��������Yr����Y+z�y1����$�S}�/��oq� ������^o�P�dء�)F����pzx��	㝝;�@�9��m�_]{_�QP=��TZ��LB�4�k���Cr,�,�QV���6�|��v/���٨��ڋ��}6��OP�_���kexjW:���J B0���
g����N�삶 5�r������&��M�)!I`�%Q@~���o5��\[$�tX�G���~%�I��V]��|��]�i#�gHq��Q4|(��g$���cA�[�ϟ�1O2�Q9����C��_q��g��~V�=h���:��ÑE�Y%�pH
���a�0��=��rM"�Lq;~���q�x��,+;iɂz��P�n��d/��\_��W>��ǽJ���R뜂��U�(���Α<�GN�c!�i��w����d��ք �5�k��E�	ѯ������_�N���m�`#q�����y�r���:`	�A�rb+��Qn���%ow��t�u�[���1�!�7�)���$��_;��A���O"�4��S�e�P��3<����FH��ؑ���lp�k.��C�Ec񌨽�&&��Ʌgl��6�1"��1t% �A'*��(�H|}Eo�-�������A(��įh�`4�<���>�u��tt����O� ���0���<��T��g�+����0I��?�<�1`�����P.J��٬�?tS����Ǘ��9�Rs��	{��QX8n��jX�_7��XP������� )��Ey���{����b�jZ~��ɣ�����)�d�Z���>�����A��(�?B|�w���$�~�db��](��P�rI_��Q�K�m��r
1*Ļ�4���":���5��;[��MH���@>���%0D|/�hC�}���1��0Y��ɿ��� �Xl-�L��G6�� X'��?����[*�G����g%�^�qJ��xx�T*fG�R|�3�z��S�(g����"Wϱ�O�(a�e�\^#i�%� �5��G&#�Ll��^�|��3<mQp��"�]���|� �~h&(�=es�{8��`�O�*G�Icn��8��ā�̫E�D�E2�D!�!d�*:W�*
���[v�0Bn�u�Kw�/�l��Kf�D-����Lh��jZE`��pD�,_�m/fF1{��ԋVY�;d�N�l�Dfw[}0��y��.�)��dP-LIo���%�b�[%_O��(�9,�lrݍ)�-�;#0��QD|��j�n,�R-��j�h�t#�?~!�y= ��%À����٤d���Wt�XѶ|O�Tp
ѧ�v�JbW&2U�2>��@j��QN��v�3���u���f	�۫]��]���pݔ����T[ڵ���A��f0eW��2�qg�~�y&dn3���ty��c��l� ܱ�� �G�W����p��l�|��Z��m����ǹlU���_&2�M��MK�XF�v�����)�y�bE�����0��l
����n���r�u6eB���٪�6�ʐ+2����bڠGD`�^���/#�-���D�٪n,Uy�3��G���6�4���c��>���,�UҀ�ј�{���+PU����%O�~%��:K"�^ v�ve��� 
fRE�����>�4[��D�J��񡀄^X[�4�[�+E��4�\rNU7F2ޕ�.K���lIT�Dnjo����6�"���&sIq�Mq-ʹΜ�̮9#���!���ɏ���׷�>$l�@_W�'��2�]rT������0�Z��n!�[�~W�.��wv�P�����2}����fS��g��̫��&��:���@ $K)�ӥ�a��u���-�U�wl�T8Dk�)��%A���F��?%
��Ֆ�v=�hcW`xL�/s���[..�����B`��@>9�LW�B�1^�[����5���|d�;┲���)p�6!�p�9��l�c��h����+v��d�=)��/�zj��a%)'|��5�1���RH�["v.ɼc�-��տ\�P�i����D=�:��6��_i�_jW��|�VU�.�O�Q�V�����q�z ��:�����E�u��v��m+��?9T��ک�LR�C�9<�u8��8���%q�!���F��M��!�_&�0���4�R�Ȃ;A���ݹ�k5c�dbw.z�Y��=��>�s+E���}�]CƢ�a�ʠs9� ��$��7�͏�2DxĢ�}aSuh���xd�
cx�Л*u���u/�\g��+Oo��yz�,l��_pV7�F��p��|����U蹋�0^ 8u��2NCQ34��k����{Ѯ�$Ы<������;�RWg��廜*�7�!�M|�\O��tȜ$�EY�p0I�'ѣ�����:$�nѵ���3O�N���y��)�l��Ep%�.�>����X$�N��Ch�|%IxS�,�;����W`�K"6\J��
G���������g2/ݛ��a��=�+���j�&�3J����&�n��d�b��2"�e�-����2�=������݂��Ge���¤-c��Q��w	;�!�)�g9=b�3����A�؍�9UL�0J�0yg������'�QIu#D�f��z t�dn�S�f�D4������Z�r�^5&L;�w,����[D�K�؛� ��ٳ������52�숝���W
�ݎ]ǧi�_����Z�p)y���*��w.g��������F�䪃0ͷ��$�yp�n)�`�/��#���B�x�=TС�+��;Q.�GmKŻ5h=�6H�	�ai��ȡ��r�	P�"]o�fȐ^�س���iȚ�/��j-"em�����4>ZƖ�i��FN���q�h�2�TtJ�O�P�3���(Z(�ʾ9����ۖ�7#���9
�h>���:���_���Ӓ�+��cF0T!����+���@��� ���7*�"�j&yR�9|f��Q~�����R���F9�d�
�/'k�q ��F�V�W�4�|s��W
�V[��1�(�ˌ���[��.�U��Ux�h���IJ+��*͕,e�!;��Q�"֗����-�	��L�lۇ���~��N��Ȗa�"
��r�B�gr�z�&��F+4�QQ�s7ћ�WC���!Ǣ��3�/1������<�#�E�x͂��UA�K���4;��j�?u�?�rqmC�����GE	F�I���e���5��S�9�W�,�sY�L�E`p���S�����[}'v9s= ��Ss���5U��t�/��\Ӱ9�
=������p���!i j5l�,�ra�>�����i豁=��J�������j����~J!F�,���A }�U��|�kW)	1^�p�����![)0���`HؙoO�{�#{��Pw��Z�[�|�����c�9���J)϶p����:T�@ 	�k�?FĤ̋�I+gr��_��*�����Y��U{�ٜ�)`Oucj5#�F)�%��0.��nd.:S�׊��f�U�g}��^8��I�x�?,��3�ݪ{�E
)�J�x���X��-�4�];��q�=x;9���`UI8 ��_(���E{D��/�{�F��g"Sҩ�����x{�Cv� �&��`b�j��i�-#7qh��ϏB�I��-��4ݗ/s�b&�lPkt���IW��S�&c�V��E�_o����/y���F��`��jt����R���=�T�'���iQ��:g�ܒ�F���퐥�`y ^����y�f�w�du貖�.)Z�,�s�*?�t����3%���n�z���K��v3�F	PHUҬSpI��kf�����!gi�$B��Ŷ��e?Ad�QQѳ�8Wm�o^=q�R���������MzI(���OTF�(�8�|�������&0�c�.�v
�4� �g՗�˕6��1�DW�/F^���1�v�Q[��ϙiD�Ý~|�A�3��}��0EeG/���S]~i�689����uj�K_\,!n���Zp�DJ}}hti906ݺ�mb{=��&H]�@^�����D�Y���<RW)�x����+$���W�V?0��'�4�*2���9�j��˚�,sS��ּ��ҖԨ�Y�Ұ�ϒ�J���m��x$��=��LW�. D9TV��G��fp��8��S:2%a3'�e��&�����t�r�R�!�٩�a�v�Ү��I�Jo��]}`�F�,n�G�bb���k -����G�9%�1b\e���D=����� ��d�
ɗ��
�g�R�eT��_��.i���p���X!�W�kk��D�>�G��H�ɠvD9�r�^�Q����i=v�{^bN3t�"fv
Z5|VT���Z��Dٓ��s�AH�&'#��l��#r��0iA�g��?��"Է�:�,U��a��B	��tc�hy6Y ��M�p��2.�o�`߄��D����_p�:�e/�-��fh+C����G�gHO�=~�<�����;���1�IlOߤ�ꁸ�|� W��M���KkZ����(�$g�7]�N�����c� '�}*��?ѱ Y�"�Ik�E�zi18���u`M-�����.��o.��l��j@�G��\b!�k��}\y�ɤ2#���e�k^����n��<�	�/`B�'�ΝK�����%��w��.��|��Ǩ�y|�D:l����Y=}d�� i��1���.�;k��� >z{�A_��s\�����S����Ww���ˏco�H����y���1��%.�#�jw�.&^�0��+d���x#�V6k|z��GF����Rlz&=/��t��.]iZ�����C�̰�2�ef2+^��b�d4�PX���w��=F��n>�z��{�,����,���aِ@ 4w�zյU��~�M��N�S�e�a2�����L��9g��.�U�Vχ(1�U ����cS�I#����`�w`6#�աt~�k�5���$�1HAp��ZN�<be#\^� Zf4���aj�]QX�Ds�-.������. h�^Mg\��Ҳ5ٮ��#K��3[n�ќ��JN[�a�G-�EUyH���
�Y�����=���#F����k�lT��
�w���7�7	*�Q19de�%���I������^x��Q����k�6�;����I������$a�J��B����w��z�$ s8�SvkL�K����j		L.��݇�;@ј��a�;�C��M��GX��qH�3�%m��1�1���zRik�h���S*u�"�2~���V�%~�!��hv�0�d��c�g��-�i���\�>�l e�o���'J�(��>���C�	�;7�9�Jb�=z�7x��M��g{2����|9��'�N*����Pt�wym�S���X�����'������0�:�U{��2m�{\#-=m��tZN˦����k�	��OV���4��J��*q�Z�bں����7��{c��:5N��uk"�P9jsۦ�h���U�&�Dَ�,�#�����8��Z�P��*�_&�����	��y��&�`��'�7�,}K��8��I��}�{�̀�Y�U�F���,��O=��G���k��G��DX7+J'�����f�]ؚ~�zl�$�R�zo!*���ҔM5�6���}�] ��v��YeQ.jV����8a6Čs�}���7��Z�U;۬-in�����������I��-���d���<[�<?>�T_���0��	">r�2@���T�E��ig��,���vŦ���q�냑�^�D7�~�b���'H>UL}��Sr-�X�|?���Y�AȣU祅S�ID��*P���� a���\[ɟ�9�o���;�;3u%�4A�f���ң;X��%��C���$g~p�(B�����Q�j1���	���}�n�c=�	�XR-x���h��J�A<)KH.M�Nق��͌h��:�$ҩ-?��-�I�+�{4e��P�ŵ�/S��e2w�YKW���1�m|KFA�e���ѵ<��F0���3��0~�mw{�F6����.����O�ʣE�Ũ��$l1V������6Bj�gY7N7���s(���Rn����ꝴt�:��:��
���Z���/W�Z(<�S��-J�Ih^zٿf�q@N��可�����Ai��]{�VW��LNŶ�~�W\�f爠��y���ƙ����g�)P:��8#m���pt��-%D�6-�5�3\�]Ƀֳy=��3�v�����qv�+���L��$諀*��ع��B���M��mhb���Ϫ�)����W��h�N�F4����~@�ۡ����4nv���W���1}/4��c�Vy���Xb��]���Z(k�Q��?0��Q[��׋L�E~���u��?���J�Z�cC�A-}����D���	��7w(�4#�麩�VW�>s�=Z���I[�GoN?�K���(�иaC��TF��]	����-��6�Q��r�r�D�F:�Q��P�û/��s�`��e%��;00�M]g��2����Dy"�M?;��\]"eV.�,g��� 4�O���G�:Bm�whf���|�;��㍯APhW Q�_n ԃ&�EI�g��H�wDe�3�I�l$XEy
i!%o���W�7ن����"Ǯ>v�XF�DN�"���C�&�jlt:S��kƒ������'M��^K��/���zz�mC���j���Z��P)���
�`�P�Ľ��Qw��}ܻ
9�̉��4��7F~�v�H5��ӻ@}(umu�1��9�M�*��l�zUq��͂����~����_�Ǽ�cΔD黼�wv����4�F�S�h��[� �/���SS���r/~����,y�H}�e����I����`6pM�%��u�D��Cg��Z~� ��p7�TR��˗s7�*���U��7��qŊ��@����C�+�AoC�ڻZ/�Y�+���j��A#,���#�؋B����z���J�.�`�ŰkF�`%���F�$�3��(�꽡!H g�ߘɮ`��&��U����2\�v��K{�����W,6���|��3_z�&D)�J�Dá�#	���寂�D�I<b������TBTA
���|���$������j����TzpY܎�:d��xD^��;p6��t�Q�B�����wD��"(��td�*s����&�����9I��m[�/{�m��9�c��ބ�WL�i����L�C'� �P�q  �ފKԅ�+"���**�(}�\_����	�.�E�b������G�QP+�%X��=l6�Q��@D�@T�I�䈏*U8��7��[M��8an��
��B��~�%�,:�'Pv w�Y���>��Q稔V�T�sQx�:uD>C�ƒ�V_�7f&��d�����-�1��"<,��Ͱ8�+���8���٪�JN��D�֭˜7PH �*�5;e���ϝ�S\��rZ9�dX'�uo���Q1n������G1~�h�g��W��7�Wo�페+�Sգv5�-�3�!���SWͣ�G�#�7w��@i�p����U�����)\KN���~�HmL��T�<Z$�>l��0�׳~�h���e��_� $U^�l��L ��>����=��=� 19�����G�_DsIz�P׋�_��[J��2W��_{rr�� �W��R:1�(zJ�v���/HL�2�]6Qs���E����P�<�-��n����:g!���� r�]
ω��V��q�3��H��~���֬F����T~�F¼����$źR(DԱf��BC��E��p��&с� �����
�����ʷ7(�(�6w��U@��>�5e=�֋-��ޢ�?`�v~6�QÛ�uc���"	ڠ�"d� �FwX$�d�7�S����}w�[�D|cQ�K�&�{<�r�h��ڸ�I�e2�eŦ���#i��EuL�(��J~ߖx�փ_V	 ���� �6ddg�D��'>����G:��25߱/�x� ��Y��c�J^��D�s}rGҎ݌-;�DѨqc��KF�S!�/�W�y�ZbExn��]9�0(���\F<T�=+<�������m�V|s�OG}��R��$�	�O�I���I5�dV�|)b���{dV��d@��;ս ގK��(�V�
�k���;N�z�f�۱$&s����.���"�<nY�A�t�BTRE��Ĩ�h�G�Z����ս��%Fm=Il�\�I�s/��r
��܊|i|}�ڤnNą�E�
b�,�X��1�p6�Q,9�rH��=@݀�^��p'K���Ş��|L�˾�EȞ��k�a �_�F�u����0a�@�{<���]�ڃ��_��R4Z�v�i(QP��T�4)�����r�y�B�j�B7[3a�5�x��d�7��1_oN��»�9�kAk~F1���^��Kt�jp�[:=�x��L ,�rl�,냯ٓ�8�̩�8�h��O'J�8G�����R# �� A��|��B�ђ1�e��>^�k?^���5E�rK�w�'���
�x>~�+��W�iT�<��>kS�?�#��/0ը��:���u�ػ���^( �l2�Ɛ�W�c~�z����B�vT3-��q#N��@�l��S�%�؝�Vpi>�
[�J�X��at�r5�v�"���f��*����O� � ��I���`P�����������8�P�߯���hR�:�/����Ă����\��f{��Sl�D��^�nv��1�_��|����Q�_��=��K6�F@�q�/�o[�>6K�#��b򊎈�[��Jd���PB�"��|��P��8�H ~�H��?�T���=�~ft�Em1Ԇ��X_O�;?��D���B/���=S��L! bw/��o��I7�?�B?j��;x&ʈ�%�	����V��}F��K7(��%���Q';����w5`�� u�e�	��K�Vw	{�&f�/'ہZ@([p�����8��<2���.����<���,N�ɽ�yC�ǐ��o�颺X���F�Ho(�$k��1]�;*.� ��<&�Z޳I���_�#r���[��m+6%Ǩ�i��K��G �̼��4��4KE�ǁ��ំ�V7wd��4��V�]��n\�Q{@�Y1�bK�Mo?V+W�p~:~��>^Y�m#aS�x^������0(�pM�xh���˿XqW�[g�ҷ�Hݜ��I�Φ鼼h�і�^�*�*3��?q]xh���T+8��l�v�؉)�E
ݫ+�,�����y�>]4���R���@&x�x�2�Y������ך����F�/�X���iG<p\rYͲ[$2��αtg|P�W��,75aq.F����*g>]ɟ�Mq�Y�Lk�,n�����tb�
'a�̖���"E��/C��ƣx�F�����ğqؒt�K�� �����0�ŪY���ƹW�܈���y������G=?UY!n�g���X_�s��F�H&��f�o��Wm�:��>(��9��8g��ط�ɣ���<��r3��u�X�7)�O��-�|;^,o��խ�|�y��}�,�d��|=���:k��稐T�C{���4-���ː�*���m���t!c5��o�Wm�3Op8杪|+�ɑ�z��}1�Sm�_��W�{�`���p��hH[��?kG'��5�s�|�u�t�6��!I( ��!Z�~ϔ8D�#th�:}m/�?��]�kY�(�xQ_�T���H��{�棅���J����|	��؎{�N6��鎁�%rr�ʋT�2^4~J�)D:o�(?��Y2L���7�S�7��Z ���z />u�0�&�^F�z�-p_ �)E��|�7)�������U�*< pю��a�=R=U23�|O�=�m�.cjՙ�+�׼�8wk?pz�UT筍��ִ�����<��#�	�mlͦ�����]�4m���0��c�O���Y,6�����m�?	{:��3�����J��Z��3�HV�w%�0�����guD�:!��W��Dh$sZ�h30�+�)D�ՂtR�P"y[�����/UwGnb��l��w>�a� ��_��K�%��3ø@��L����27�"!٤�;��g$�
,3��k�n��@�'��ge|C��~�Z�!@�.*;�L81��!{�z.�(��[�Tq7 e2��qG�9���Ƌ=���e�_�@��I��}��u�+���(q�a_��b��J�h��'\�6��?z���={�db5&�7
<M7�=�'�IY�E��<��(oRzl��Q���]=�%��M$i�5o�t5�Qd��5v�WgB�!D�����.�$�'��Mdv�K*�*lC�c�C����z�����}m���F�ʃ��	(��uö�[�Ò�-��e#�k�]�J+�ߖ�45�� �O�f8�T<�8�1��@��-�KdUl�x�}�.Pz�,2\��DŲ����MD�>��Z�������=�>N�$���L��Q�����_�����rb�*_
뤦ly�9���x�NOh���H���{��KQ���}�^���ǔ��,	���Ậ��?y�g���(��y�ZP�K�+��o����$�cԅ�纝�zMәxB��-p�UB�KXC�^��H�iv�@�`�w�kM�N��4�&I�\5�fD�9�����d��^I�6�od�ɖg�/�'�Z����4�����(�ܯ�.�z�7YV�}���O�/��.��b�Gg�K����kݦ���o(^�!�vr5YA����}���
Kp����>o����11�8IN��"�0*��Gx�@~+u��
��_�^7OP�I�&�:�7K�Ӵ�1EY�$��2r�  �I���{��*ӇǼ�sRY��˕u����PbU�h��� �,WZ�С��\c6��ѕ�-���4 �f�߷�C���1� �<�wܘʹ���y<پ�]�+�L����^��;/^a?��H�:F-ԋ܋!2��bf�'��1��e�����Av���q�H7��<�( Q����R��^�c��OV���1v\}+� 4pr;�erӚ
-�&���:'ݠ��1�~�v	L�P8d�fĒUE&Q��Ƣ1����tCqRt)@#
��gR2o�p����<[{����N8	б2���M���O9�O��p�>�".�a���D��s�]em�d���a?qd]�TՐ~&�N�4y�Ӵq$�뉫6�Xу�Mf�y��x!Gת��l�����E0�$.��ӫ��y���}cGݑ�0����(���?�
f�:�����fV�"F�3+:�����Qϧ�ۤ�nʗ����Ƙ�~�ώ�L�'f�p��	��>l-ڃ�!=|�!���M���Y��ֲ�;y�6�'��2�3���4��S�(�}T:q�-�d+�J?���F�s��+��w��z��&��e
狞4* ;�h��H� 0�Y�bT9ཌྷ���YWq�~r��l�����(|)2Dk�&dq�|���3��m|u)L���K �ï_n�g�J�ߩ��( 2 �R�8���� �)';���
�h���rk3�����`�X%�hA*_L�m���R~���#�+��as�/!�orx��p�O<�;���+f����o���N#������ɤr!���"����c�v-�r�0wG5+ߛ�mt
M�^J�H];�OeeǾ���\����gZ�u���!0��.(�h��{%��
�E���k:��r�дZ���r{x�ƯI"��E�-Y�4�H��鬃�%��^6�5&�L~��G\b���rm�B�r@�	�)/��q>I�d���rGJ�w<�̿��/Z�X��ʍ/�2eټ�`U���
+Ғo�ѫn���O9��d��4;)�m^7���?�N(��Q}f|SF�5R�����:��?���e�xYT��q҅��#�w��2OSN�T1��f�92�n)eԡ����z��ś'�l�?<�) a�h� �R3;"�vs�[}'�L��>
;T���`��i����n8L{�OUu$�J����^PKΚ(t�Wvқ;�3����
�fvف���e��z&���U������d�T#����K7�i�BY��U���Ӏv�YV���@4�a�əV�:Z=E��T�b�gUDzN5�~�D:��S!1�H��g[�uPS&��I�7�d�#_�I5�	�X�π]�=���RQ�i���k�u���$���/�|��:�r4����^7Э��HtfB�7�'�J����%<�+9(���I�vNH��󾹤�`�j��ٽE�%�}��r�x����9��_�P���a�@-�\��R��]s����\��8c�9ݱ�Q����D��U"S�Di�(�p�t�#�]�?W���xq�����ŏ�ܩ-�!b ��E������'���X.�~��u�״�QA����E�XsT���/��Ϙ�";T��bYG�y�]Rf,ۍ��r���@�m�_�Q`W�PAo6��gb�!����-o�Ҁw�f���}�'Yc/<� �^!-`�$+��í���$.�e�踬���\�N%����IRv1��t��"�#W����!�K=�9��
�P�Fj��P�P#X@~��r���C�7x��P+Z������I[�y�G,�ɣ����Z�<���2!�pO�7T�ɏ,�m��N��C{[�D�vY��N��͇�3�p�*k����ȥX�Ҝ���#A�G��ML'��I#i�`��b �U=tV��0���9�B7��g7h|����ҫlB��Z}pX�Q�"���%�4�����47.�q���m��>@U�!�N�>^A⦕��lII�/�g,�/���[܃�TRo��	5{ �t����˞FV/��k9��/���S9g}��!�F��p�ܩ�5-�NԬ�����N�����g���#x߄�-�Vd�@���?�%#�A�`���	�->y�	~��9%�&cM�Q��	`�����f�OU92����g�~y���*�e���c΃y>Qyc��O����f.�zW5�]��8c7�{~hmBD�<ͷW��"6�z7�+5��~&L�г�b�I(��s�Y��7:j8�c^Ok��%��w����L{���F8� ��
�K�2�W(�l�n��0W+q�����׫���f������րi"�8Wk���V�Hٶ��u1�~�?ХiF)������v���C��V�K�1���@ڻw�<}T~���(��:o�����F7����~�^�Q�7e�d����@���j:(����^C�\�k�?���eB��-�SFk�̈́�6��t�[�����)Z�����N0��Z���;Ӗ#4�ây
~��`y�V��"ig�7gzk,D��z��:؝��'��u�v�唙���t\Y'-u;�e�Xݖ��Y,�+�R�I�j$����_s�CQ�����=9�0���b*;?Eh���������P�($��,1�����pϣ��>d^��u�WY*�IX�Lɹ�Q*��F�LyH&�
s;�R�T?��`��[ժ��d;.v�4��Es�̲���R�}T�l'E�#�qnl^�`8��1,��Q�F:�Ё�1����h�v�6]�+q%�P��dj�8�u�|5UOjyiCub]�%�b3������V�����ƻ�&6!�ʝ[R��0�<����"�k�5������t�!��݋X+�Ꙓ����,�0,D���;�δ-�ם�օD�2�1'_�W�����I���^S����&!i�&�o^(D�*M�Yō������ￖ���l�������,h;��@<��G����s��,�H2u$Q�-�:/`�� ׊9�{�%��:�8/��mVD��N0m%7pV��82�X兩Z#K��?�GR"N��akڇ#���K3RH�򛸹pm!ys~�?�jw	�4�s�d���
�_/ �'�#	��#�o��5U�IZ�\S]M��y2�\3$�CzV5{*����ŶgK�*MԮ��)��!�Ϭb�$W���a�'��� 5]�-8��?G�7.߾�q��<w6��e�6�  횕-$�G�Hf�¦�_���.��!�K��8�6[۸�����gr�}�_.,�������S2�(?p���`[�t(����jh�K�gPٓ����=��dB������wȫ�6��eԹV�`�.�:RI��y��0���aZH�S>hD9�g��~a}��i��Q'f���ڠu(��e..�R@�A����KVm�*�|3�� {��ӿ�a}6VJ1��k-�j��V�����M��S��%^&�EN�Pj���q��A/�pK2��;n�1IO��f#�A��N�3 ���_㥢�w�yL�љ$�G3�	�37�r(N�~�ty	>{��{�J�,f��e�^P��%Eg�ԋ+��^���Sob۬���.'4-�D����fP����V��N�q�[pS�Ǔ���t�e���v�G���c]&���8EX�h�X��[��cu��*��z	rF"���������ȃ���^�n�=�2�+�&_�9�|Ԭ�30�-m��WA�:}"�����*q^,K�V���Bj�u2����fxI�t�	S�� �Y;K,_�''i>���
�%`���z�Ag��c���}��bQ{�y��h,o=}H#H,���/��^W�dmEatB.� 񻝎����'��3�[�f�z�yrٜН1&6�mŲ�f"�P8�w�1 ��t.�
7�Zl����5E��kԋ�N�^7��n�,���]*�ܷ�U��{������("��v���%�%���k��n���M��~��\���:x=��}�զ&Uy&�Մ=�R����8>���4�k.O�cq�7k��חR'����6"܅�r�6 �B�P���
��ϴ�����E�7=�"3�V���@y���aA����埏.���MQVE�/S���_�حַ�*7$�f�=s�U��� ^81%�J��p�c��{�/��ȡ+��N6J��V'��f9��K�{�6�Mx�O�Qum[~\sa;����݌{�c��9�}&?���ma�lggݲY�F⒵�>��������}fc�^<��#�{0���OC�%a=\�o��ڱ?qQW���u��:!�[��~μ[��)�H� 4�@<�0�ݷ"
�)~g4�h��H7 ?����;�K��,�������
�Jd��+�/� �i�x;�׍���9�NA�̷3���GD�L����q�g`oH���a0��&_�&}+J���<lBaE�J��F*���m;Q�"����vn㨪|�.��󎺢�,(t T�!��9���`ϸbno�5�uǮ~*e]���ز�m=�kN�c�'P��)x05݀kWr�+���"�!7i+�8ʐ�<�eV���$�U]�d�O��@g{���R�>G?��`Q����36�z+���G^7,t�C��!85U�a��?�[@dsz��F''����hKP�{ ؊_$������e�!i�w�?ٚ-�mVg�4�G���K���=��ܤ�;�Bq֎�x\�z��m=��V���ʜ6�"��%��j+r�G�k��.��9�)㪔4���	�N�[J�	f�Z	��1��������|�_�y&�rp����܉5����0��tw�wÆ2��:�%c{�ޗ���gQ��D��b�>C�^]�}�6%�ׯ�zZ���mj�L�5%e+�6��Ԙ5��ݖj�A��K�a<CΙ4�Ǽʪb 7Jf�E�ƺ��}x�;��_~a��.hx���5�S�ۼNɠt����q8p�U�.D��~�'Ђ�y��F��ݽ��xa{'�������[�Zr��	���9P�pA]���Wlv[\i��}�ŉ�z+������T�;��㔗����2ܤt��G�'w,��T)�Fk=I�7�0���[�$GV��a�4��Kˁo�s�����_�0o侁>�k�E���eٵ�[Uy��tI��,+�.�m�p�c��^��/���	)��6�G{�;�r	Bq��{�����=����t� V<EC"��e2�ؔ�p_eT�
�A��Ue.%d4�U"�Sޕ'6z�D���2u&6�?���RS�se#LKV��2GA��ѭ�'�9ۍǆ���变�`�R��s�}�(,7ą�������޳�����֘~���
��Y�3O�4'0��Z �r'zb"�q]�c��۬��Z�-���4+��"��t��8�oU��͎�N��ǃdGb�t�o;��XmIhb:���u�Y.AF�J�����oгbd��?> 8��ْ/�po�?�zVO��5��`�M�D�&ۇ��m������|Ȅ���wMN���IkBz&p��^�H,:J溯<O��Zr����j�}U��eO���������}���ʲ�pX�wR�˼��et.-��f��cy�hB;Hc"T�P�*�-��qT5N�$ǳݨM3��ƘaWu%��^�E��J/��Z�5_��n�33Bh�?��$��;V䫣n��jX��qyj���!��z��R�/���w?&��m�lc�T@¥T$�vR��G�{�Ï�_�`�iD��T"����x
nGؑ��S'*<%����f���{&{@4"�m���q���ߋ�/��,e��Y���6b��6y^�Ke�{�%,��zW#0�#aC4W��i�0�7W%*H�J�Rč��N�;`6}��}\7�R��l�ul�L{�y�j�`���"���|�4v������)���ӶU�@����I�a9 ��N����o�M�ᡭ�) O�t�Ū����q�9˒�hR��b�i�*a*�wôn������`�_��Qi�rH Q94����xv���\/M���+�<w;� MY�Ũ�.Z�T^(d�|�$&���{��B�*"xw��;pR(�ʁ�A����k]�X�~ S�<��W�p����CZoH��5&����=0n�b���Ι�w�	��X�f/������Ǳ
y����������b��}*����lb"����>�����D�f���"r��P�Mg����|{ޓ��u�ˢ;"Vmj��y��[�'���[�o�]���?�K:-���N� �p�D�k�Jw��K��ՉXT�>����	AQ�(���ܴ�	��Ȫ�q-Xu�3]庣a3t0v�f�օưfGXA�tj0�H]��	����U���^'���.�r�2b�P��!�$�ݩ��PXO�a���sn��AN�[���J�3��ێu6��2��y3*|'�s�M��̂sߕa��I�@=g���
�S}�?Y��`x�?�tWݫ�A�<�qL����BPٗY�x2{N ��5��;5�@os7��>�F�%�/����RU%�)|��&W�>�xC���Ċ�f$>:�.FO�1K��s7�c�|�h�̀\Ћ���kp�{�Rѐ_�?+�!n�`: �v\�޼���4jD�]B��ҫ������[<%��D���&�e�A;{Є���� VH���������tkn(����%���ڙ-�a�V�|�x	=�{B�o}�	����|V��@h�������
i��&,�^kmC��@W�"�ɓ�0���E�������7���g�}�z�>��e6�{X�z�#�X�K�s(���<��L,$���Pv�Uv��1k�m�յi5G�*6Q<og��ހ�a�;/�Z�#�؃�5̝L�9 )��=\V��D��(��]�u_��N9����G��2UY��Z6i��~�P���x��l߬_�w�dn�Tv�Mc���<�4ܦ$������i�s�d���U�9:[�s��ՊA� F$�ƴ�?���O�j�����N�߿p�RH������?�=��#V`f�������E��7J�l����%m }�z�GIQ���#.��Ȃƍ�7Ɉ�9i��00���T1�����/~�\�	�M�}���^�׆{�B:ᰶ�]a5`p=��r��c�S�jeC�;9&;#���{���QqM*��鰢�N����q@���Ƌ��@vq���oы���̮�绥mҳ���]���J�u���!Ԏ���Mc$�&������@,�u��h��� A��4�fx�C�G�D#����a�u��i%+��]�b`Y���&/��c���9��w�MGQ�~s_�϶��ͮ[��Y�� )��W�S���Ծmٻ �P%I���ݜ��[���h�
�Ly�7����m�N��M��%��YB+��n�zY�7vE�!	W��"��Y'� �L�d,c�3	��nk�T��2��[ ���X;4��-m�� 鲛����{\�yԤP��	���
vj�;���~�����V�ҋ��
��R��fcP�����0�e�����|��+Y��D�w�UO��ڐ��R(u����@n�%%܌�%0��:v���������A�͸�w�M�&��[�uy������qu���Lf��@ ��vG�����Z�J���l��Y=u�[�x֙0C��i�<�ӟ%n[��w	���Lm�
j���Ż��� ���X:o�>�c��s7��ȎrҭM��M��V^q�������M%���l�8Tp�l����<JZ�vz�����$44ĎUQ��O$�������*�hO_xhW1�X�l���e��,F��&���\��1�Qz�6@�j]���>9�^�}��tӑ���tD7�����K�����ra�}$�k�����a�i�g��gV��X�<L�'l�����N���O	SO'�3�o��55�ԢI$i�T��꒥�
�U�Oo��5p�2��"<��]h�J�\p�w���Scʠ���l�S_n�h#>��EA��,F�n���vZ��P�e�jG"��L�n�s�^)AW�V��	V��1�~��Wd��&k�l4�K"�4�/V9}"s�v����\Ehy����evs�%��v���y�0�:pB)��K�Ҝ �Z�@ڳo���1|j8Z�yc2� ���I�ڟ�R�.��w	���l�@*�?�{9�~���@��0��[i4	����EV}�zy�,�Y[��<r'��r���}A�3��wXYT�M�ߥ.�|>l���o1z1�8 Jd��vX}\�~��WgD�/^��%����dN�nk�3���iƘ� ��Ͼ5fkc�B1��(ӣH ���Jr̽?����&| y���-%�G��!͊�)�+�A��p��Y�s�p�9<�X����_T(siW���VY;��U��E�`h:p�#T
aOںE����Yʍ握S�<d�d�p31�R�(������������JQ�xyzu�m�$�.~�[���Ė�8�� ��j�/�*^&�?W��+�ų�8M-v$
�}��q���R�t���xW��cA�*���V�wC個���Z�J����mz1'�"X����JLRf������U����\d��5Iu�nMZ�V\q�D�l����'g���
!�� �
�����j��Ag�
��D�G�xt�a2n	��^�x�7b� �n���n�4[���֯`�0'߻��S�����R�+�gq�.�Z�"����߅d�,�]P�>�x�y?,u[&�$�)p7�x��Q�f����f[�M�b:��$���2�V�-H����`B V�K�qC�42�? GJ���v����I�S�}��@��G:���h{p���fз	l��߃���$x/�O_w�%	J�,e��L6(?=v�}s1L�s�:hl��%�rc�#��M�E��k%��UV�������	�f�E��3���*1NW]`NQ�/�>�
qި�������4�-��,�,X�N���M�m�\O$�����Q�dQ1�������U4A��7��d0�{i��3^YU�t���e��W���=[˴��IJ�����_��f���d���y�c.��B�Km�4����ȓjH�Y@e�j����'��L���M�p�?;¿�'�9�j˲	��4nN�ы�ݾ̙����د�t�Z@�>��&����ˆݒt�^��	���ۆ,�aj��-�9�}D��A��.�������qc�
;v���+���e�ƴ�C�B�\�:�G1�:��F݉�ºl�Y����§�F2��j��À�8�>$6thڃ_
͞z�sPy��v]s��F�)�n�E�}]�U|'�k��XXgE�g%(9����:nD�}m�o��7ב�WM=�R�i 	��� `f�u�M��J�fY��@��n #,����Q���`�H0�(��&s��~����RQ��5�oY&��>})G�ϩ&����L��E��}��Ue�)�Η7�S��<���n|�b������<^J����aV����7΀=���9����ʤ|��<i'�ܢ��x��V��Zz��Ib� p����D�Ԉ Q̡�BP�lL�
ώ&Me���M�U��~.��D�'�GVe�?��_���ٷ�`0�G�ֈ�i^z�,��KT8�f<�.
QYAFxR�X�'�(/q,���2;�m\�|Hÿ���*!��d!������^Y��
ɴ<_p�K�g��1�֥j�O�̀?�0�8ՇC㙴@���U�m|�*�h��C$AC��;6�N��ޢ#y�0+Ƀ���D�U����Bᚹ"��a5�3����K4��b���!Olv�>��U|)����|5�v�~�8\�����'����L��Y@�o^"��锚I7���N��-,[����6n;4���Ba���O5M���
�[��7C��AD�灍�L��z��0xJ���-���dAT���B��I�3�I)C:�TQ��~�=Z�˩f���-�:�T����J�p��ݾ�^$T��ɫ ��G���C�n@g2G	���r�|�pz�=�/�>o���)����7��e����4�a�N0� �|�b �g\����ڶ0~�P
`_�ں�|�ێ*&��޺�����Ш��N�I����d*�9]�ݒkW�T�d����<�j��TP�(9�D㭥Bx�F�2f��Ŷ���LS�`���#E<ĴK#&ʯ|q����W���m��ajjꠂ/�K�۩�" ���'S�S���:CL��0;���M�6"�@4�s���$d��-$����n�-"��t{�vf{�c����$�YA��Ѥ����d�*�C��)���/�.��^̘�&��Q9I�F%�������'�-�}'#�ZfFeý�-�2ݣ��X�o�=�?��]\��GA�. �X��X7��5b�)����e:6�*�)�ď��{��"��s�r0�:ּ��w�yL=e�i ǐ��p�܏em4V��U���p	q�wqIy���i�Ye��3��{ٴ�d���n(*MR9&�����c�x����N��D �0�E;�>d�A��g�9�k��)��Uu�i�vQ�?ʸ#�X*��_��F~��N�-��!���~��s8�@}�H��$y��@�hd��A�m�nI�2��19��W7V�6��"�Pg�ϻW�~���lX��:Q*qÝ�j�7�S��Z#�ұ���h�N�З���m�Wk�� I��WiL3t�����P]^������塳�6�m�1��6��2?9f��c��?}�E�N8�e�!%,��B5�m+q2�q�Z\%׋�4��������\r��ݴ�[@�h����*�}�At�����k����ǹ����y����� 5���E&�ز���:P�*vrl��Y�S	��o}7����6b���_o��U��D��ᚏ)���3o�>t�U�J�}d�h�ʃ����Ƹ��[��|���v|k�X��i�{&:e̶�C"D+�#��k*#��i����%l�h�5�G{pj''iV-�1ZE6�\u�
k\��\�&Jr,/�o��o�$�-<=GtR+	�(1o�;67G����kD�#1����+1C2��_He(c˻$�9U} m�����Qv��uL���߫JU(�/���~�_>5�O,MATZ�Ԋկ�V@���ă�`��Ww,�������i?�('�N���ڀ�O�b,^�5	���^5�Q��<F:.YĲ�������w	���sh��
��p��H �������f�������n��p���M閱� ���`X,�^:6<9H��	�=,��n�S��f�VA�4����+�>8@���8x�������>ï�N�D�P�=#���|O��Р|38�V���r�,�Y�s�6���߰���ئ��kAW�������;
]���Ç�d����G�TuIK+�Km�u�w5l嘓�2n?~���˺����3ؾ/}0\ز�U�^�9/��-~�}�o�
ɮ7�X(���:�_��߹�R�����,B+�S�5-��B�HF���ŵ/��&��"^/uL�ڐd 'ԉ�#f{��>(#9���-��"�Λ��M]J��~� �w3��vV�[~ҧ���g2��0w���P��( ��6�����6�4�І�ph=�`���a1αQ���xVRȑ�0�&ŵ��<+;�S���0M�$���%�`�;�s5�%����MSle�4��R=i���\Jf��_@2[�~N�n�W�����ݐ	T2�&�'�M��us�U3Vv�b�;��\�� �m� �|�ScJ�D�� ���Y,��1����L߳v�,�0�˚�f���A:Tw<�}^��_��F�>껇@�
oʝ�Bu�0f\f�����__���c_��'~��,�+�Հ]FOl��a4��y���o4�֢+:$A	K��u6_�һm��5E]Ѷ�1�:L���k��������`��˞Dq�$��<���Jo�|
�m��i�@�j�4t
G,�%*<�<H���	����,�y��[�hv3I٦��Е����Y����K1��c�g[����P�pb7U"�{��_���;�1	���(2���Xͭ�0���m�'�Hc��C �{��:k�qkl7�SN�8 �%��^�4y�{i��꘯���]�j��D����U�wFR��mji����{3q̉8@�|�c��T��
�̅9�݈a!''pnѓ���T������vV2�x��b\*Exm�,?!�p��lN:c�3��$��(U���'I�:�g�#����S�b�T��?�)�5���'D"�1�-�HĎ��0I��(�N�q/tӑk�Xisax����A���u���mi|c�Z 4$zrsr;he������YE�J�R7�!ﰶR��t�`G3�C$r'.�,P�x:١�������dY�8�ZTQ��O �>ZB���<t���W�ݕ�u�º��?Lyɗz��|Au�$h7��ɥu��e�P��q��}�ሗ����A��ds����M�����igv�_Y�x���L�K%��6�,�^���7N�u����]����Ӆِ��gW��O�������zn�Gy`��Ѫ�S<ҙ���$���ufm���֠!�&`�q�z�b����؝�����p�3�R��MӴ2�$��x���x� �w�\�F���pl�gAzE4�ő@�qʆJ�\��*��t93�w��� �In}��������P~v��nh������`jj�̫B�=E��;3s��T�]�;� "�v�mv�3��ү�����U;b�ߐ�ٻ��5�vj��]~C�HEZ4�kq�¤zc�@mr���+\��[��QC�:8?���$v���©"�@��ұq�[���H�u�T�b��,8��ۿ��oȜD�\4�������<�^<�0e�IT��g���֌��L,��sGn/`���t��}�� �� ;���8Û��Y)H1w��&�QWms�怦*� ������P����,V��6G8��Rjsm��*e�i �y7��9����Y������	���LӺ�k��^�p���?.�P����j�N�5�=Y�<Qɾ�ε�ㄿ�o�#����sŎ5�I��xM�7�^�"U�g�g8��/�'���T�o����f�C"������P�7�%_�x�C99cÓq�����H���,"�9�:���{�Ai�o�� ����D~����%�+U�27u`c��Qvl&|��6~�S�ڸ�AL��"U �����iA4���9Wf�G=D��-��/:\��%�R��e`�q�St�%$��ր�	��T�`��-V?���K;7gI��%�j�1P�V�QCZj_-x�?�>�tT~��-քC<jj��9O��\��!�ȉ�L|�8�IBX��*J E��}hj���l�^Nw�]�#�狃�U�i84|Tn�)J���YD�5�����K6�>������{�ЂC��V7^X2R7,��KQJ�8"�!)xn��x�4��B�;�HhLI�DX��&	��D�'�◰X�.�q��'cB|�N�����fjw1\rmE�o��>5�X{|yH�'
�j��y�-�0��%@.ai�Zr1��O0�+�K�^���V�dޤ,q���I��344҈�p��4��M�A���ο�3�g�`���I��j@OA:��ҟ�8�p��=zؖ?Ո�?��z�xyl�]�����xB��c��"4���5����v��ۅj�'����u���+��n>�=�R����'Mp4A9=�]���EP�mx��$���p��Թ���Y�<?�zTcW!��Lz����#�J�@<Bg5Q|�+֞��q�4;�dmԙ������Q!�U>�	��U<���HF��w�)��10_��ZGj�C�8ÏOkl�u�3))���+��Ҙ�D�"N����L�5�n�����(�!����,��9üL\��(�r�٢oʍa{���滢�pT�ۏMU���;�n��Y߁��_d�A���J�WaN Ңv���[ù"�U�^4��Ĭ��v���
��b���wn�]�RAτ6Kc]�u��!*&�b�0n\�v��q�*�ha��_,M֙�aJ��k���T\5�q���0<շIng����7�����s�9�$�L�2��_�k�HI#��)�<*Mռ��ˊY��pFB�A%��8z��F�x�Xȡ�V�ޱ���0��(H�`~��/?�	�����$���:��r�>�Oj�D��C�/ڊ���d�]��y9���([.f`��s�HjH�����=:5���Z���e��y��D`��S���!�@�Zwx�9�T��+���
 �4$�� ��p$�)�y�H������=O
��GL�H>�Uy��Ό�z;�3�&���xUt�;VX5?�@t��H`=�	4�rE��<����U(�%�{�>҅ue_OF�S��k�#me�k���%+��u2h�����iR��q&���ٟ0YK3٠�� ��E�ڸ\䪪����~L@�_.٧��&ܘz�����*XcKtw��%�o�	p<�z)�`?6gs���F�\��!Gw���X��g�x�/I����1稰��Ν���u����U�O�%��^�g&�q�M�"B�mph�� Ad�*��s��� �B�	�YSGU'Q�04�����o�IU���,xAȄ �S�TާY׾RH�t��i�� QsX])aPBw�%�V�A�V����Z!ޫ��r�0&z"�M�8 Ñ#�i��`���̀oF�����мN$�8���+i�*��s�����
�c�ù:�xwT՝0��%�37�ͱ휍�h��.��yW���@�]��~���f�;$����}	����A�e�W�oA� � �ޘ�]\�X;��\d��&W�{��X�;��1�M�p,�=�d*�~H��~T�n���B���P�j%0-�A�4�!<���]���ܰO�V�K[Ѱn-Sfg$�왷�*9IJ*���H�4��uy����Az�ɇ��U�#��j�9�d$����S]_��0���UTE]��l�|��P-ȉq�R��'V�c���-SI:Bg�rX�{ i;�-J�N��s�ݎG�.p������,��"���D�'�d�`_N�u�ڱ
;K����Q"<4������Ju������rTG@R�Z�5[���0l#}�e�V������t�i�@B	 �˷��3��g�Z��q�f-��cl9��`�{�����]/���1Ѱ��O�GJs`��"�A�,����v�Xե'���Z���sVA?/��R:-�#4��	v\m^�-�5;�9��]�Y4�l���*�j��E�O!l��
�r�Ӎ"�l��>q7A��E�)�Gا����2����Ovq/�h"�%�q�3p-�X'	�'��%�-G�P���ε�K�^�b6��vM����\ز?;�Ȥ==���
��{8��:>�h�]��u�&f �8c���a^��T�sF�k�4����F��$�K�5���Otwl������᥷H\l�_�y�$�)�ԃ��4p]!&��|��ϗ �("�ۢ��hdͮ�����]���+֌p�g�z��^��aLrAۅ)�Z��w��zTx(^��U�o���cx���y2N.�P�j25Z�_�5��H{Y���A"�霁K|M�fkO�K�Y��_i��m}��鯵�sJ��{�����9���r:��~�ʓ<��/[���}$	Ơ�ڬ��)PN�B���=��G?��ٮq3��#e��y�j�B�U��"~ٺD!���U������\�!�-e�!�@�k��a�/f
D�K��`S���(<�q�"7�p�mDD~��y����b�����e���%�#'}�T�P��fԇ\�9��صJ��P�K�˺0���X'��7�0v.�x�f���\dJz��K�����|,N�o��L���<�-�˫�t&�����oE��ap��
�(e���/�	�客�Ҷ��=o�����{�~=�k��/�]'+�]$"
#gF�k��h؏����$����#���ܒ�>��Ih��fDf@%)�RX'��IF�`��:���X�������OqS�EQ]��=�n���������O}:��u�<^}ھn��x�����Ӄ̢��tm�n����'����O~�.���i�ّ?Τ�n`�xDUp�P'�T���M�(�瞉��B���\�X˟�Ib��ۃ
�M�W�i��,�E	yA3�	��'��yB{i���Z��
���{ilT#���w/V�lq/���f�MO��p�2��r�2A���e�dR�a�n����h�R�3�bW#i�����/Ew�54K�@�k01p�WΨ['
X�Ӹ����}�d���U��,YO��?)�P�\ �:� 
mg�U����Y�]2Ln�&�e��n�Y�a#�L�3�|�n�8�#�����V{E���OC���b����R�����Ӗ�hvt�Bw� ὕ �p�j9�@)�*W�g��CL�������9{��?�\,��R�����|T~�L�ϋ�r�}j�C���Ӎlyv�@�L3|�[����ܕ�W~��M�R�F�<�=��Ȓ���E����p%!���C�FU���t�qAי	R�����+��5ٲ��J+�i����j9i3�S���
D��C�8����L7~/8|Lg�.*�����%&���	tz���v�쇹 r���#���A ���I͢�����t��;�榙�>�t�kj܃��u���	���@#V�'!��)ѻ��Gu�j�R�"���{h[��W��w�v��(�k��B��b�Ɗ�ă����Zg��M���]�
E�qZF;-{��C��#>ʚ��K@����k����SLnR�8�����j��V��b�B����=�:G|Q�����3���3�o��{��"�v����C۾2�g]ŉ��0�;�Ò�+�/tK��]�O�������[b���l��-#�xF�#�c���k������:�o����i'hZ�|�����Q�'�E_j�i+�j��]b����m'@#�7�$
��:)�q����{5��#��N,�����������@*c�������hn_bb��
�$�G�Ͱ;���\9��kF�2W�3��f�y_WEk	|\yV�@B��耻��6�#�
 -|KiYXw��TVLZlb�=yR�~�j���#^��&����*b�4�Yy�/^��b|�i���/�-���p��V�xpW�ͺ�^x�_��A���]�&�(kz �����Lq���`!�_���ׁ�F�T����9�ic$���z�xZ���� Ƌ�9hm\��LX��*�,DaF�'����3(�J Gux�g~��_Di��iV�I[����>~c�O�q�o��Fӹx���=j���*�b �fI�r+�%LY"=���P��jH��}�V�B����]> �2�;�Į��V4_ؙ,��lJ}��{���p���5X{4(�w�'N-�	�DA�w��?�Xs��j�鲴���ȮT�l-�N��qWcx���U���<О�	�6��'�����{R���y�m��?�]�f��c�K[��Y].9s�8�.L�����u�IO^PU!@_���K��������b�@�_9m6��� ;#}���oK��˻H�Ml��Q���ࢺ�p5=N|`��a�qjp�ҵ7��u`��%�=���[�d{���M̥���6�}�y}��\�'d�检چ5��!�Ӂ72!�/�7�J�(ɒ�v�Y%�����Q���ea~�t-���u ߼f��'a[u�'�A[-5�C�x��ty�T] ��.)a��I����.ʄ��g� �$�Q��2���k���p�a.�z}��"�����5&��˸Y�B�'�i�V���D*H�RA)�se�V��4ZВ�99������1��H9&Y�u���؅vr2P�C�W����W��*���);]i�Ok������[�F%;ש���o�|�^�2f3%A���H_��������:F�z������CH�f��<�~H�k�]�&��R��^T����ce��i��wN� ����w��"�2�/�Kz(k��{^`�4��Ɉ\ZB�T���[�:�ք�,㪜��d�	��[tp�>���"������fFt8�P��q��;e�4}}��[��K��(�b�]̃�y�][���{��?����Mp�*�[6������2Q�J"�Ci����-b�e]���%�[ ���?�O�zA�H8�j�����y z����B��q���݄?FU���*1H�M�{;$	����-f�����?S��!��3���pn�kE��PDK�*���b��P�.��Fe��nc�G��3j�N��i��Ndl�ć�^p�yA5�T���u������o�5��+�祩{��� Du4�-=D;A4
�U\�J�w����C�=��e�ڛ��?�HKS��`�o��Z:���>X��%�@��ӊxU��YP,{%���q 9ϱ��Ø����jT��ٲ)���t��]�y�I�ޕ�
Un7\
�\�Vk�U��+��Wl���#hM^ǌ�J�	��ICA*1���uM)W�5�]Q!��t	�p�h,W}�ή����	�\�=�w��o)�G�Nh�l������~���zj�e	�'�` �jՠ�L���%�nFJ*�>�^_�!D��fIW�<~����1���k3E(�$m2I�1�	`]�Uiq` g/ O�g�!R>��O�z�����;,2��	���I�م���uz&,�{(g�"��"���9��h���6�����2pr�ݪR��3�U��%o+�P���h�@����CG�q��=�=��EbsثFbl;އ����m�������R����,~�@��:Kp8C��85P�o�����w��D�������1B?�|3��!1�hr���>׍�����pAY�;Ȣ5fkjFه��X�-�f��"C\��W¢�b|{���z
ZF�Jy� 0�2����D�L�u=P�����x�Ѝ�<�C՞'X}�(p�׬��X�t䦡5̍�ö�פM�D�`-1�8zV��2�V�`��F��+�υ�Ӹ��2u�G��P\�b��v�Z��v��DG�G"0�A�Z���@?��4�bߊ�D��[���Y�Z�ghZ4�.�����TT����Y�bDӁ�zwp�I�����r�I[m�%t�F�|O�=�5�H�8����m���}�ސ�q!ܑ���6̈��������7C~҈�@�|1s���q\8�� aj�9a�3F�RE�Fh#�F��������g+YQh�״������Q."_���$���P0z�Y�����k�-)�]|LP����=�*+��z�s$T&�i�|� N
�Y�e���1��d�P�u:Gre��S���K]�F�
�N!�U<�g�w�;�ђ"��n���UlUR�
�G�2���"�k�X�3(�*ӈ�OASfr�!9y���r��m���|zۖ�� ^1
�ŮX�W�u|XY�Е�[�.r}����7j���+�r�#Z�2�5�ԯ��=Y?�3 ��z��W�)
�~�����?���Oy�������C&��`�BB!��,\c�@��NX�1�|���\�����i2�B�ƈo9t/7m��̾2
JW��J$��/�u��n6(%^�:
���SaN>���e �1O�)�f?�v�e;��j��<��"�Ұ<2L�ɣ��:i��N>�q��j<��<���4�ŒlNW�=e�sY-��o�x��	�9&0��p�YE���ș�u��6�?^vI/��[��rn�j8f@��k��H\6\�b���_q۸���ń�i�����8'��\疤R�kL.�e�m��c�	�I�\��}��h�ׄ�N
����fа��P�ًh�+�����5�H#����ê@HNl|`S�! ����=c3���1���F���rp����X�+��b�_�М�FsFA@7����#)�b���J����ٮ�e��Kd��pC>>B��,���\�� �]��O�:���P����x��r�릜��O̭�����ަ�)�@V�a�O1B��8��{�[�-%ٿP�e9z�Κ\V:6x
���;|�k���8[5W Y��#��i�f�J����	�����ʹX;�j���@H®+�?�A4�<B��qJ_���S
2G���T��ZnG����j�{%8J� F�I�w`�x�9�<���2�`_CA{�P��&l�,��1l�:T�>m��*�x�TV6l�5^��YtW�L�2U��b�� A��ER��QE���#�����?���+S�k��I�L�'��/ՃfW�'%g+4t	�������� ����<��\,�w%�ue�@�.�=�!��\T��cс���ئ��c��uC��2��jMl��82���q��}Ôd�3&������D�+����|�Z���%��f�����R�B�����6�wuj���Q��D �I;�����{�}���í=�|+s抄~���$�]Xl��ԞHdؔ�I�^(7w�ʜ��0�e�����0+P��^��Neے"'������E���9���`����:�m7.AhV݇ץD��ڄX�9�황� N�L�P!`�'�U�R�)̓%b	��ㇳJ�
����<!�����F�}�fo�4e$��Du�e�X�y��I�闘�<��(��*)y18-_�5���ڽK�~����©�$�'�]�"��`��<Oȵ��e�>�z�XǢ�Q^���>� 	%w��	�/��ċ����I8L��6u���?���gp��{T[�)��&;}O��$�4�7I���?:9�d��VO>fN�Z$���`
�x�(3'W4]N����>�Z%r��ty}@��E�����xV0�
���a$<R�K���&Q���Գ"&,k���p�?�JD*�$v��V�y��|.����6�@�O�$]K�X��ˁ�S��\b;��T�%��iIki�3�\�	�wC�����4�M�&�$���\��`5iCr�R1n���:K
���` %���3S�
H�ooP�����
��y���k�~Km���֙��	) ��9������m�0E��v��Nʃ�V��:Q^51������������%z; 
������k�ь�O�3�
�q�[]@��{����{{�j]����#�-���h�'AG���*^96��B�.ߨ�/PD�'ܮ9�;V�5�yl�4�
:K4�Q��a�Ԯ���:-b����}/��B��5Xm�ʆ���Ţt:���KF<���(o��U���9b �҆��z����'������'p�M�R��<�2C��N��'��p�3c��2��gԜ���0v�t��-a�n)�L�c�0�t9n��V�4�}�A��=��D%����z�3�h|�Y�������i��8G)��ɴM��ԗ�IE�X�a��囯z���a�G����.~7��
1�{�XD�ΕHd�`	=��"�u&��!Y���~��=��T=#W\k�o����m���~ī���|�L��G���Ʃ�#^� ���T�:�HS�6'%�G�ud��?ܧ��*���i7�ͦ��ˢ?��8���|�k�a����F��A�v��$&u��cm1���L�郑T�,�Z95s��\=�I-c|P@��v��<��X0���h$�#D��djۣ���J~fH���(�7��s���=�=�ś���̩ږK�X21���M���H�S#逐������6����ep��5w���G�H��b�^F�|nOASUx�lc7�����[[�<�p��B���A���}�6T�+W�q7I�)Z"ԙ��k�3��{��y]��D�D:���	D�g �1�a��4|>z8�u \�t��ѩ��Cr]��~d�쾣U�J�1��G���I�JW�>?~wnfӼb��:l��d�.�a���B�-�d�/(t��ݙv������Oഽ�)���a��_�U'i�׊wC/�H4#��Г3N.M�H�ם*��5K'����t58���ڑN�/��o���R����CWj�d���|q�����!mEUmTm����R���tc7+I��,p������9�^h4n��N��Ԭ��$d��J��Pl
��p�dz_0_�n� ?�� ��_nw�ee8�z-�g�^j�y���ݗߋ\c<�߆	n|�����v�\�����}��ϓ#�X ��q�xV�3и$�ŧ�`�U���,P9��D=bx��.YL+��fw�$OSUE�V*v�������\��}D��d')�I%�SBx�xd|���Ka��
\n	�QZ�P�Z(,-il�E\"iѽ�l�����/��x="Id]�ά\�d���)��^!�ڷ�ј�֣G�������Ղc+�p6�Ɵ��	u�����KF�î^�������*�J[��������)���+N���7.3�۰�����	�l��o\C�����g�4Q���#Y�e3��)�GM���� ��s�}���2wڝ�N�v��I�G�	��hoYR���--C�7����M�u��L�ᲀo0���%�V,a��/|�)���d���ol���ȧe�'��%����h�tɑ���M@�AI@�94L�i��0,٦J�&��@ƎN�Ǧ�P��~/���O��H7���^s`i��o���f��M%�޺3Jz}��S|��o�oW��wǷ�����J�Q>�E�'@����=�6��֥���{��,8j�j�+�r����iʪʺ�jYb��ĭD�˯B����d��m��v&c��M��*�O��~�%\(bWh@�zatjm�6�"�7Ru�R����;���T�h���gWW�|r�:���,�mo���������X��G�Z�[B-ґ�Q��@��Q��tc �V�,�@6M���4�&�L~��a���������Ѹ�q@���\�#x�������$쀁]��&h6|��aw�>���E�v&��Í);��U� ��*&},w,�- W�4��Yf��RC�Q����(�
�Xڗ�[	m�E^�"�9� ��Z]��)`���6#T;���O}�S�b�ݼ�@l��b]��Ń���ƸEf��)L�uY�Dk�[0�U:�~]K�~�L@֑�١�Jn��8���:X4�%��8�fJ���`�R%׷��k������,8�5���qӞ|�#D�k�{���i��K�g�uD<�?������P.	��x-&� ʆ��J��!]�: ��,�I4?և@��4:|���Ξ�o�8H�^��K��1�yU��f�tQ�RH�Ε{v]��>;����:�V9�PyΛ}�nh��1�uȔ�,��7،�/^��v��ïk�ԎEIM�Ȣ�]����	@�ήʡ-��U���u��2m����9�:�^�sK7�|CQ��(F�%�4<np�>�8 �/GgN(9_I��p������j��1�9���Sj�#��f����/���l5$��#Z��?א��[�9a�KиO?�u���'i�������G�]Z�wC�����0��(�¶�5�[�κ�xQ2e���+KI d��\7x�T�$r/���Ӏ�����-���J��JC��rd����J��O�����"��r�ЂK@zu�@���b؋lX��A���pp���X�.�=���P���|)�݋^(vs5����g��'4��+]�ҽ��f�6]`�b�ږ��,|��p�Z;$sAV5kF��BGL#w�%5p�Et�m�,]%�ELu�TYv�}ך���UJs>�	d&u*�����	-m��3�K��@��$�s��٠WRN�f�x$��s��"�Q���������7��~�|�[m��`A�GCd=GK�o}��ɼ��r�H	�F�@<a��&}0ܭg�	H2����ٔ�S��o-,M�vKF��D-���h�z����a�zK�%�6�β��)�^��b˕�A�����c�����2�`#)�0�V��o0�hj9נ�W�&���{�cG�2���f�z@�v1��)2@�f^��0�wn�H�Z��Ҷ:�y��B��D%:kQݐ|�(���t3
��F��XyHT�I�{;j��9Eh<�u���4�%z�\� dyU��j>4�#-�������&q⏰�m���,���Ȋ�7�LG�_�`�����2�F����0����4[��w�
�8gT�^K�뚁�69Ձ���V���#��S��#����i]N�v�J�>�Jh�C��Q����}]+�����8=Mt*Qg��]���}���u+aͦ�"?�@���q�Ԅ��JH�A�,�.q��7�,����^a��ox�n�Yos1�(A�)Ã���0�sn�[O��"@{�}��K���H=���ɉb(Ƈ������*4[��'b��km�c�6^4t�Yy�����|�n���>�8C�|K��v��^�g�^{�|d��f6���F^B��ب��,���g�W��7�%���J���#^r��`5I�9���$�w�"�=�U����ŝG�p�&�G�';�H�nT5�h
x���3F�������nU���iEv����~���'Dvx�c�#�"��)|�=�?i� �����t..�q
��8�R���Q]�]![3��I�	���,H۶O���(�����ة[`�����:����Q�����=#A�w��Q ��'Tr�m��h*Z����z�4�!���H�/23=��Q��:���A��j-�kM�d�m�!?fɛw3�3�Lw=��Ү$;�p������s e�p��͖�(�kw�e,������ԁ��.��M�u׊m,)��[1���f,�]ly>̞��a�)Y�r�#ǞԼ��
��#� �.~t���Z[@���1вY-���j>UG!�������&ķD��C����z0:p�Xi�Bsig��?��ըķg�俀��Hg�S��)����m?b��sGm��t �0�㒻�#�(ڦZ �h���s)�6&��傏.y�Y�ɺ�L����Vk��(9�Z�ΩP��t t�q����Y;���_��0�Y��:rh�ɫ���	�Ɛ�v�`�c��R��v��B\G���m;�`��h$d���i�P�)��yi�/Ywg8H�b;� Z(�5��Z�5������ڎ��LZ�����ƶ��Ff<(������?ek���߁��4�.-�b:��Z��=��۱&���G�^��ǋd3�(�~V�%V�8C�AKC��]M2	�ު��%`'t���+JQ$��]aT/x #��Zn�9�uQ�inJ,>�^�SB��`����a�$�����#Y������� GK�uIb�:��_7��ȑ�Z(�*iX	�Ļk8YrY�,oLl<v�xXv�������r��HjZ�̳+r�������E(�)�m�Xz�5:e����[^�Op�-c����ηu_6'[Зy	����3#�"�l���"���]�b��9Dp~�/;7��N+���rt8�.\H\v:�+U�kݐ([�i1dV��ɟɐ¦l|k��f��Qɉ���Q�
sK����f\�ˑsʾ����i�}����`�d!���atn*��4�#E�9�
5�yo�t���~]�I#��oĻ��L�5F�^�߇ie���Q22��e2�Q%5*ܮ�t	\��`��.�F��]+S!ۨ~�(2Ǭ��0\�� �C�����XAeK.l�_tԆ���U=ρJul*%�D�ɡ�:�Ɯ3�+���:W��|_~3�,��s[�w��!��L������bf!0�O��MdKj�ǉی;��n;E*�^cW��9�h
�h!h	�m�q~�4��ĨP�/��M/���H�@E:(2�1�w:~�p25�]�}bf[�1��_�] ?�ﺯ��?��Z�<a��-�ĢZ��e�1�2���X-4_mSk��KV+��?��I�Fߺ�����~_����C)���i!sޔ+�t�u�0�Ɠ��b��?y��T�D,V�*���@E��g4�M>�]g����F'3���"����а�����k(�G��2d`XOԿsա�~���O�P� ݬ�&�-Z`���	df
E�/G�����s�0���������=nPh�<�bA"��p|� �� ��"G��N	���P��������^4MpF��6~Lՠ��P�H��wix�s�߀c����px�Fl����N��$���o<{k|s��[S���s�����2�ш��÷���\Ojݩ�j��9G�dҀh���	��\��WJ����akCe��������?��D����\N���ttz�/�p?3��»(><jQӛ6b�w��q�[�ݘ����@qB@������W�r7��W��:��!�����C=�r[C�{ye�tKǽ�j|��M��?t�޷�4�AQB�!�;휎�F6PTc�� 3M�$�N��4������P����s�}�ա�O�<~�J�E�ٱ��V�GX輼�y��7 ����\��r`
��/�N�&�_]��R�)��E���A�R9(W��6��Q��9��J�A��*�2L�"����m�J��)��*��G�$bpv�HɵR}�����g5*u)���N-�0	&o!9cCGD�%�|��|n�5�����W�(��'��=9<��Ol}�(���-Lhj�=��ފ�a��A\����Ugܿ>�LPZ�N��5Ր\X �a�W��p����I!V�l�����G��En Rp��b-Jd�hlM�H5</]�|���n�dp(M�4m�g3���g�hQ�f�g�@<�����CZ��Y��d�Xj���>æ����0���Y��<���\�Oz�)XCn�cVM���ο���1l���t���L����(�{��e�1:ɮ
+Y�?�ewU�F�H6ʒ(a���[<x(y�1b��3�q�O�78
�&l��(��Z�dP \��ST���B
��J6kC�Y�ſ*�23=E���!����?�
���(�C.U�6�3�����)"��Y���ē[@�Bݿ�|���m<x*p�� �_��Ĝj2���or�5˘Y1!O!7)����/-���$���'�����1��;˞���IU��e��R�G�E@�Z���B!Oi+��8�e2v�op�5�{�N�4.|qdL�	� ���P�l@��`Kv���X��5��),Đ=�1ծp4V���}x���=�`Z�ıdP�5��u�vJ�^�y((���؝���֑��:��������%Jм��.�Z�).$����ZЊ��Y��x���p��Lu)��u� n8R�E���lZ�=�����\qa�|˺p~�
t�][,B&�Ї�~Ƣ�]m'9)E
3��[��f��W'��E�����­Iy��`�8ءة���U��fנ6��l{Ï���I�˧����Ȋ~>\���=��9�o�c����M4����9YD�q��q�p׏���E���}�%Ɏ�Q#.��N)Ƭ@]Q���;.{���_wz�K��hsxh���z��-fk�a�θp�{�s��dږ5��TUIؽ~�gv���_5�!�\����ڎ���`��3&�s�1�
��$[4Ʋn �4������!q���d��qۄs�D��Qiti_�uv�C�Ē�#JI %cc����h8���%���-�
$��N��Zz7�!؄�Y�����ű.�۽Ƽ�HɅ� �
�ʑQv�"��Qz�W�Q�
����~������'pC�@�̗�%���=�Ei��s/q��:�9�&c�7�ԥb�4��z���rq���l=�H�v���EE	4xc�r���`C"�*�e�m�񽽪r1*P�Ӭq���a���DF��#�����QBs���$�3�U��7ۙ��z����F���Q�R�K"��_�7N/����k]%�K&YՃ�_�]-(Y%z';@��m#Ȇ�sm����o	�����?�ԛ Jr	�{�֒ý]4TBVu (u���_��g��ԁ�Z��C�%�fX]�����jȌ����5��Fj֡b�������U���+TW2�j�;|�:�����*`��V!g�Y�a��@|�q�;�FN�8wX�}8���L�Q�	���T�e��H����*h~�4U/A�}��o5�Ui}���A�[y��`���*GQ�GO�w���"��Ծ����]e�>���@�� ����d�*��~�H�1�iuۨ	%�&�x����W�L����T)����'�iP�@�lj��`��.�`���%������֥b�t��������=�,-�&@ �٨ߤs�@I:�Z͇�4"}OA�ϒ���f���@0Wq��Zaa�1��ȹ���l����q��szɊcf�Bw��r�["��u�P�	��"w1q����u���3��*��z:����:�b?	mю�x3��z��L�]�8��E�s��k;��Wϥ��E�%��}t���`4�_%�is�2k�8S'�$�����H�\��m`���1."�v>z���=�����k=ZԤ�j��~��SQ�=����G��.G:�pGq�;8|k
���|U"L5f�Y�ˆ���P�]DH�+�|�^�w�!l�Dhl}��s�����K	6p*�+�;�-Mn���{G]!�2m�͚�2!��ː�嵙�1������;��7~����B}#8�^O��6	a-
��q�N����GPJS�׼7h���*��|2�[x�"��n$�V�0��Ͳ�e<S-��S4�l�U�K2.4+��	Ȗ0���5�N}x��2o��x��(���>� �W���:p�e�W��a\�jI0�.Q/;8�/�d�C����#���66�@*���
k�hG^M�eD�cw�i\�P0X����O�'7$��1�1���/��-ʉ�uM2�C
�!t�^�J����u�]��!ܓL�v'���������U����Y8�̮�N_7b���_�~"�R/$>�e��5�Q}�`�7�@мK �yis��Wh��0F(8ֿ1��FF�M�,[�ۊ�T�4�p�42���X�&F0oG�/���q�L"T��!'4���i}���
iZ�wO�B��f���f��������4Z�z	�%�2=n�k�~�pE[&�z0�4�~=�h�dh��#���\)����6V?{�Q]S-^i1�T�����'멛�[ѣvաLݏ����\�@��yM�PY���p�+�[�
�
����&��`:O-�������.K�1��(��D��c�\��4�B0�1�-�c!7SD-���F��L�*��c����*O[�=�c&���]�~l�M�#�6a��o�����wp?�wW��=F]��[MF��[���4`�HFH(��h��Du�?�8�d��zߗ`O�Ƴ¿���pf��u���M��H_o�C�Z�8��k6�� )t���m�I*�6��8md\ƍ?���̭��H^梕�f�jq�D�r+�Cy5y�k��Ak�^֔n�����B{�	7(�u`�:���v�p<�}���R�R�]yk�
|M"0L�����6�S�s�Eݱ{����|�XS>\U��s9a� ���\�������9:<d�Y��.	>Cۖ��N>���eu���+��@���<>U$Yj��P�`:�6ZA�G���}>��"�-f�糱q��t�p���0cb�ہ~K�1���
g
��*ȷ��]������4�˕yrq��`��M�\:�\�/%��ؿ����G�i4�D=�/I�m~^���4�z�?��õ��k!v�����QBl�Lf���_'�w�d-�ҩ' ?/�����RTa�~	K:��S��(�o]��u�����q=�U&ut�ox�t�7�i�U��~/���.�K��f+O�.��n����5�(O�Bk߅�CW�I�έ��&��3Z#�:)3��PY��:b��2[��p���L;�m�c�	Q�0�x]�YT.��2v2�6�k��%�_�
/2��#`�)�H�1yڌ��d���'ŀi��X0��Y$�R
s�~~���7�o�K� b!M�~Y�Ζqr�ڰ	�5[1W��u�f��Y���8������Y7�!�Ϣ}�5a%� �ƠA3����=U�V��y�<L�#�O}��9=3�p�l]�$��1.5�I8wA���W���X�dխ����c>F���z��{j7${0A�2_�	��PQ���Ә!XB�3%co$q�$����dӂ��x�Z��${Ģ�ILv�,w��C���X^-�T��3�D�̨���5��S*��ʠz�fL�%���)J����
C,��OHB��y诏^��$��
A[����V{��#V�s��"9*�0�W��4	LUAhmK�v7�<�g:���J���7�f��F�9F�����]��\i]�&i��L��� |��(jϕz�/4>tSH�#��㘅��;���ѻ'AR�؄Bh͗zv����P�6�,Y��k&�	F�Zr~q}�L���W ��k!�Xy���W��-McӣHB�ѧ�h%�T�������OB;Ud:G�8M��s�[dg�"�Q�֯���B��ټ�%,��M⋨��8��]	����O2�7���XN��#��;�u�Lc����I���*Q�3�ߍ=]����z��Mm�i?(>�܏�P�[b}�8zރ��S[��s����&�ԍSs$�X�H0�`s��թ�a��Z�p�0b%fJ��c`S�06f�f�nW���������_�����U��)�yǽ/�h�"�5$����Fܐ19�E�La���u�1�/!6�r9�^�{�$ٳ�v��y~�[���P��s��yK���I4�;��3�|�/*�s�t�^Ѷ�4�k�Y;?8����
T9J��}:��T�����w��g��zS���s��ś��*{˛�'����׮�����n	������㯵ݶ%:i7!����q���hV�D*ݭ���a�9	nҨ�o��0-��4~�a�'iV8 tA���*l�������}��ߊ�S���E�Q�75��*%�=�9qӽo���� �(�#G�������9�ٻR�j��yk�������ϴ��P�-JL����r��n�~�#�������H�	�X=��>��ֹ����doD�H����G��#>����߲�?��bV��c`b�&��W�˨C���������WV�@������9�����a�
#\��:?s��� ^h((���؃�Y�gaC�V��	��-��l�/�Z	}g^i�ݼ1�!�J�3�q;>����ɠ��ŀُr��MFӸ%Q|R!J�!L�䎽�E/�Pq���(��J*���T�� P&�����Eէ	��@�5=cG4���0;�m��V#U��_^�%fF*�dUI՗\Q}Ioqw��4-�g4a��	ٶALsIk�薽��+ѷ{���5�s]���^���r�*��H�Nw7�'���'�JOtW���L�u�I��6�^�g�j01c\? |����@7�V�]��X��k�ѣ�ǝ�͹�dLƪԮ�p};�:_Z�|$�2T�۞QP�V�$͸d�Tv|�����$R(�IS4�=ӳL��Z�D��M!Ef�l �Wq�-a����3Gdnuږ�64S}���l�y��m�Xt]�le
�0��#�b��a[?��9���b� ���@%Pׅ=o!	�s@$L�F��yGen%
O������4�ڼ.⊱�t�<|ۀ��y��Z�R`�|�ltp�Z��,�|�B�d����r���Y�8_�	�F]�� K>}m�K"}}�.f`���W ���ќ#Nb� �(P�а�2�ORx���b����'݄E��=ڽ2Y��~�U������V`�SF�<+�c�4�^ˢ���Nn�<]F���� �>ChF�	����� �3�
�� m�(�,�@����ꏼ�ۢ��Rj"�]�z��k���آ��R��~iq,�q��S��d|"�AjX���.e����zJ�%���z��N�,em'ԥ�_��g��Ta|��T���aIۘ�gݯ����ن���V	ר0/��9�X�y�Ux&�Y��Krk
[Ŭ��~�Slԣ)FaR���<a�����6m))@M� 1��h0�^o�s[̎�r����@<�bK=�K-�}��ܝ<n �߅l�NL2�i���t_ʋ���^�qډ�r ���u"� �!�h��~r"�{	�Ȝz����UX���d��
�2�{~=n�dH�<D��7��D܂�9�Uv��\3-n�z�I��<�����䓀G��,֛�W;�D�8_�*r��em96H������>�Ēw�X��G�$�;�<�
�M\@J8O��u��q<H0hCG^�w}���愖���*���y@�D���,�?Dx��(͍�Ӹ�:s��hٞH'%j�BkI|"�N�%�&�hX�׿��l]�׀�[��0�Fw�eW����}5��w�
�� ߟ���M(wcO��ϻ��W��sͼ%3��S��/#���J�!r��������P��x�e�<�<����1� �c�ژ�ǥnE������jBߞeӷ��>�VdEj5���oxx�&�]����({�7:�n��2�a�@��n��"��/��+����g<�ܤÅ���
�0-�ʽmζ?ƹ�h�]��7��%�R�ZM���TOd�"��Z&*��NU�0��)���E�������,���~?Q�c��L��ڊIH�q�'j��[�&����Si�������T\���/EU�cM�֛���"�'�J2����$�5^����#q�H�T
�a��Ǥ)�Wdu�� s�Ҿ~���{e@R�s�8W*{�Z�l��	˜�0��B�����]�6�oی8��mCAqN�\Wi\����Qs��ɶ�_R��j��4!�*������{L9�J�sT`<A����PP�%�˗��K���k��qA��S
��K�I��g��|���C�;B��3N`/٧C�%餩���"�)�~V��- 6���{B�«J, =��	;�q������Q8�LX{վH��d)��&
4�a�}z�~[+�prF��RW���9o8̱�{����\e�`��#�0.˸T#��Ί5z(�=@���?�;&�@�p�4�3)���5��΃AĦ�V0�-�ݟ���	�2�[1�0|�p,��F�m�)�)�!I�g��ۧ�$7N���^HW�����f������,�O���������?.����9�.�*{��g��"Ts�4٘���N���������U�G�.�+��+�=D:����?��>:��}_5q�/�?.��UM��#��6nҎd��eD(��
�-e�)���ڥ�����������M#�W��E,s� /���D]�?.}hb�_[��r��|-1�B�͕��*���u�u���m�> 0��4
=lw�>�6��hy���Aq_��\1���6�z�V�Ya�'5f�5��N��Ah�Y�Ǖ��u����Ҕ��Ă��z�r�u�ps0�m7F�eѓ3��T �Uw9�F;$�g���<sg/�nJն���%s��Y���W�w��~�ߟ���v�[�hT���j��T��������߬��D���T��D��E�a��܈$C�g�J�0�c�d�,~�=:�p�@~��=[�عG��Mz��J�)󸺮i|�1Ax���`�/f�<�+�s�����eY-Y/�rY���G�}g��DO��]}�!I0�ZTAL��iX��F<�Չ��f���)�Ŋ��"r_�@�
�H_�IH�"�K]�(����C���k����k��Y�O�n!p���A�'�ZH~�Üm9��Z��[>�mB�M逤v���3�Q���,����-�nZa( ���}����3�^A�����9�y�%�/�:�UMs���\>z<´؇o���gvp�8���g ƪuH�9��>uW�gO�^�qb�z��!���g���D>�{�)��eײAD�D��ռ�m�K^Gd�7( �Nf�,��őCw!z0�����R�
������� |�;g��@u�9����r�I��/{��+������������ŵ7_X�ܔ<Ck��p$�@�����"�z��/ 
#�o�0�a ��}�?)��ּ4T_�jr��FA���#5ï��;Zn���Q�L��:u�.G�$7�'�NÈ�C�ŏ���S ��5ޢD����ЍE	M8f�+�B��&!r9�<�m��,/���P��u��Zͫ�t�m'��f�f�5��N�V��Pt�%,����hbXQ�g�ӓlj�����&��pԻ�nǒ�ї�_���s�-Yb�Z8� yWg�R�<��f{�C͍16�D�1�^�Ӎ�tֱ��Vvo�Y�*/�����Gv��1i�+b��U�$�󷾹���+(������gN�u�!��-x>D5�,��"��$h��m�n�)C��J8p��'�jE�w+k��1ZF9~GD:�t��,�N�Am�<���K�75��@k� K-1[����	��I2Ax�����Q��ă�cm[�S1���^�T�Z���g��*��t���>�o��6ʴ���+H����*ꑒk�:�>�;9X��ۣ�b}�RJx�βä�#�0C��ߧiu'�G�"�-9س��`��'��eP�����寃���)(X����9�[�,���
��X���+P^��z�<����8������Z�����w3��$�cE�ك�t-{�I���[�bF�Qf�MT+D�t\�}ȍv�6.��Vp�G��h����j��:eZ蔋؈C��Q�"QQ8��8����V5�o\5����b�0��\R�O�J��T|�����'�`#�w��No(�����B�j�Ј���~����N��4�n3�����"z�Ug'>�PǁY_�x�i�=�Z[��fJ��e�����rZS�-�`*��_�������oo5����%����:�e��"Su�#@�Ã6����o���ҷƸ���?���e�}��#��>
��;�詷�K�y��@>g.�U�������/�o!Uhsz&��>����p�\-z��Bm�d��#���Q*��bؐy�CU��⃭�������}UY�L"ί1ȿt����y�

�j�|�y��0xJ�D�6#)�7�B�A�HC9����iz*�NsE��qٙ�q�hbq��~�dQ��ml����>۩v���t��k��.�^;C��2��$Şf�#o!�.�s�xp˅��Y�|tl��4M��Mn�t���`����-�#6mU.N�ɀ�'q����p6�qc���н���z�@" �fm���#$�?_]�
0Q+���]G�"e�3=���P��m�r\F�y�x�9�F���{ԍ�#L{���~�:����j�8�%S�j�][���<�54�}�e*�ne2i (#F����b.2�s��J���x-	��4��|�*:�<6����E �=���Ұw�R�9�0-�	���$R	n1�.{�G����X0\qRʐ��Q��3�u�A/��?�ov}: 7J?��6�Ms��՚Bp�sh��/0i��*_Y��564
�6 !��̞i��r8Ǵ��8|v������y�D�l�kz�B��}��e�
\������S|jQ$@���h�C|ޛ����S�n�E�kq[�`P}Z��aRٳ���NbMrA�
��{"VhkM���6�!�(��޾C:앏�;��;�S>�(�@y�lЃ����OdQ��h����[K�^-:��!�dT��]*�'��.��՜���s�H-���=��QJZ�1ޅqZ�y�K��kT{&y�>^@t�R������Ew���z~̿b�E�B��=�W c�ȫ�6̒T^J�G�	c��G%�>B<�B��6����ϯ����(CDx�����n��aY�B~�	��O��H�.A��l���9�1��fH���L�a:t�f��"{��TP_�,�C�F�3��?��{XGIg5Е��)�i�oǣ@��$��?�|�7M)�s%��*���~���X�z�~%����S�sL����P~hl�dKsED�|\U��~ti���h?2
�_�	<o��tK��V~*��P��0x?*|�ю)��Pf{I�ۋ����Vs�,}�0C����U���l�MY�&F>	�x�VF9��\n�\�%�V�.�y�.�ZB�)6��Rf�I��ˉ`�8��e�S:�eGQk���A������\�B���=�?���Y��Lb�N}z���=ɞ�	v��+��{��"&�k�l(�6��:��_Ǯf%^`y�VZ�l��v���-'��E�.�^=�7%fP�cC�*r��\��A��qZ�$�431"�Ԯ��?a��Iat���!ab��Ƙĺ��ە,��[�c��!��������G����	����� $\3"���:y�*U���K�4�M�ǐC��l�H�?�6��P��{���"�.��Gu�EƹE�����@���Ǥ�	�$���\(ڟ�,���(Edbis�?"3� �O{ ��,���[P�S��M�ȳ���5��B�s�Lz�Sm{��o�z�O�:i�XX�ة_�E�g�M�,��,�u�0�ٟ����?a��xQf�!�1���B/S���Dtϟ1G-��<��-K��
�=Kv[I@ƿ]$h=b�8��X�L���tv�F����5�ŀ@�8S������_+�h���Ĉ���V*�Ad�`���UK��cR>I���R�'S;Vw��6��_>��p�@�d�x�t����zc+|=�A�G.�����4�6����S����q��Fm�������镕TP(͖�`�}�'ij���}�h�w���5k����G>��s��2(��9�t�፺p)"�A��mHei����MD���:���bʗ��F�a�oJu%�Ki��=k��������v:��1�\0�\[p��E��4���W��f��]u����Э�yzK�Q�ǣar[���AvC�D��2�B���Ύ��.V�<j+������>_�hPN�`a�;�4vM6�-Y
<�k��Jy�E�?��%U�b�<5|k��[���K����u>��������������|�o,���ME��I��Wq\O�t���]y��l�,q��]C�<�!�u�3�i�Y��R�n�����Y���/^�
�!����v�B�i��|�;jVQ6%�οv���ݻI��P�C}����'U�:�v�ѵg�p�إ$bV���f���@߹�iN�'�7��	R�k�Ǚ(�Rbp(���D��O0)9\ЍN�c}��~�"+��vB��GO��Ɏ:�67������ߒo��FBs�󮒫%��:� ��!�Կ�fTXv�^;t��-��T�z�ѹ��mD�v/�E�b^7 $�.����Sx'η�N�ޒ
��@�ԓm�4�KC���a��e��d0���%m3�"�M�A�0��X<}�gJ�L�q��pݪ|��-����e��o�C�K��@M��y�6��J���}�
��W����s��fnb�$sE�*�Hf��(���"=/I�\��R����g�o]`=iBT�E?D/��h�)�c��3 �/��@���ǒ�������ɥ_a�`�J��w�UD��@��5&I?^ӕ����T��/�H����H@�k�ji}$h�\Y��)c�,�>"۞��Ӑ���Hƌ�$������V2w0S�h�#��D�8���2�m�OZF�sx~y�^��A�%�������e$<�պ�'��4{�
~��<����\'؜i\�]I�2�Ԓ�����c�9�s;��%���md�Ȃ�*MU^����2�F&���ρl���*���o�`c�!\��Y�4�����|t"�ȍ������ ����q��Ғ���y�h��s��F�HL/H�� �x�U�y�p�4=
'�[ׇڣ�#�f�]�.4*l��	Q�oqٛ�� ��Pn���Q��*�8C���vPi/p6��>��tӗ[omf���lߺr@�|1�/��%�~�	% C��xsp>D����Yz2�SF�w��¯DsB�F���uЮ���qR[%�k< ���Ӣӫ_��EA�0��v���OƖ`t�Oq|�?��L3�z���z��&����������9/������	+�d@@F�w��W@�m�'�H�;���?'(��\�#�'"���͓xm6vpX���1�;R��p� HX�p!k�\\^�ZJ^~�?�o��Ne�?�M\%�z	v��V�S��,���|S��(�ep��22	.�:�?`2H��]��~��g�%��ȁ������ҟ����*g�9OPd2�d<%��4A���P������jHm�`���q�Ύ��e�M��Mj#�͟��S�-�s^�H�ZF��C?>:��3n�^�f}%fd��ڃ��B�m��h���hH� cB=�Ԑvה�eh�+mOm�~�cj����PCD�=`�:-PJ�"��i�v����&c�'r����E"{�y����"r'� =X�,����"B�g��2�Y��BǾY8�/�O-���������z�A���z�H�.�!PgS�(d�&x�&�$�X|�B5�h�;I�c�Ϝ�w0�o� �HH��*%�Td@*,g�]�Z��P�5��$��aC����W���#gT=f\û��{W�D�� '���ƕ=�&1.sɢ��L�q-P`�~���<+��P�	�t� ^����m�*Ӫ��L�X=�׼�f7�퐲�|�xU�C���B�ӵ��e�K�8a�2Vfe�O�6��ɢ@#�UM�n-N�h�.���?�u�~?G�����y�bO�;QR�|�i�Iҡ�o!�(�����p��p뇅�hf���_�W�/%����C�BB�;0������ ��;Z�k��7t�75A~�uRj]B�u���P rD���(y��a�H�(��w��.�@�d���(��~	.{?-"�& 6e"U��o�*��!���^�BޢG��$&ݧ���-Xu�'�R����yU�4����ķ���U+�-����HP����/�LA��E5e��pt.EC튬}Q~�`^�i&��|+�!D�4|ci�W(x风<�.����k4X.���IP��E�2�&"���AE��q��d;)��?�A-q�����f�fY�BXm� I�;��8M��ϋ��̮�@I��j*5�.�(�ʨS�.[c�W'�z�ߛH������Â�[d�,@L�U�7.D=�)o����|�x��5޹�S�p?��+�.C�p�N�G"��bn����S\����k�@��y�����X{F��O��]�T��e�5�Lh�� ˳�Lmv~�ɹ���M�P(��t�Z��G�;4��wUMfWпt+�:י_��tZa���z������6��/b�'��4�"IH�A�λu0�*R*j�N�+=h_x�4ٞ>��sK���.��1yM��d�V��U-?l{@�V-�#�*A��h��9��xfPN���)����wd���S�CKa��x>��*\h`�g6�D6�b���¬�ҹe�w�B$�*Aٴ�L���72ҵz�7���*W�����U�U�E�Y�.moCW;�����O�ôaZO�����(zb�����&���*Rnw�*3�����AVp<���E]�j��;���]�i�v��iV[�)F�D�+�5s-��ڸ�|H󦱼�����`?aJ�Yb�=R���OjGA��Q��l�݂��y���4�"�n��a<Ӊ�3S����r�6[T��+���EMK'v�n`�}�� l��s�;̥Cj6O9���|���#^ū���� ��F��I1P6Q���)������kj���Ot�&E���S}�d��ZE�G���j�1�>�E����Ճ�,G�(�;��Y�Q��5��Rj#�ڹ�\_�A���i	1 e�Ul�
����?r�6���wJ�b(��v����錐ۆX���k*24��]�[V�����0��[0P�z���s(]��l��6���Z�����Q�=Ą���o!�#����㋉[�qK�"#�pDz�����"i�f�5�z�`��.���J��<�K	��#���ȴ�n��7&|��Y���)~�y�Ժ^b�=j�HުG��N j�m`y�w��4^��:	TQe��χ�����;?��`w��ҀZ\��Ll�_�Z����H�w�h����JE��V���䢌�E~�S������{�wo�I�H�(�K�:�	w��>�A�8!Ә�e���A�2dW��s�J�~2�F8 q�YH�.��Hp8��i�JlD6��'>OtT=��)�qAm�L��O�����
L]�l�d|������)p�Q��,['�TK���9���ʟǨ���=�i_��͵Kz��F`�+G�:ݘ�^1�F�p��v~�8��*3Z��җ�un/� V��a��u���K��Y9ά������a�ܗN$�
s=/���> ߴ?�ĉ��:P���eB�XQ��؊�$Z��s�/:zHU2`���	���I���W<ŝÒ]��є#��y���=��e���s�U����,��1ʉ>	�姸��0L�ٻ�o|D��ҋe]o3Xp�����_93c%�AQC;�5�o1u'�"��~����D*�J�	[��Sw�X�uN��!��vH���lר�]j������,�v�에r��D\���+�Z�[%k�����j��g�� ��K�;�'�{���I�s��+��0���_|�$�@؇G��Е�r���"jw�r�� � ���D�h�Z��ǚ����6f�"dj�ҝ�Z�!�9/�V.zٸY�5�TRf�W���=8Fc��A,�ѿ��h��H�<����$�#F��Յ��<t=�w�"��]��S�YRԗ���@-H�`�n��Zo���r�ۓ�d�=Q��vs�f�5��{�긥?��]���]�~�;v�m�,��|v4d!��y� �L�G�clN�a��]���9N�=PF=50¸����+�iq^m�Ya��*<΀�������;e[�2iX��om2�$_w,=����u��j�C����(��Q�u]�>%�v��u;�����ñ	Z����Jk�J3��8���Bf�$;�T4S�q����n�G��u�Mԣߵ�����D馍`�Ѝq�_^��V:�"4SW�>��g�tD6f��=S|ΓC�ܩb�`�m�kJ83�w���������V1�2m	b,h� ����A�H��� q����l"�V$@��{�u6[�%�n8���2�ޯ�Y� �n�$1�3���7�Qj�D��z�H �k���Uv|D?_uu��<�j�%�͛�E\1Dg���ь��� �:o��h��CP+�L�vZ�,6��LB*��A�]��:D;���}�0]���0(��H��
D�BR�EPPHJW�eC\��9.;q(��)򍴸SI��\��ݔNY�;I��7'AAÄǫ���b�e��-%�ad�Ten<�����+;��Z�'<2J�f�_�b��[�[��{��4�zY}�<�Z�a\X>�oW�k��h��I?�q�hybI$�(,�Z>�	Å�p�K	�!�!s����T�{��a�o� ��-����1C:S�c����$�l���b,�<��+y�= ��`��a�o��q�9w�#��ܽw�L"j��n	�C.��В:���m�G�g�[�M9rF�I�cB�^������t��%޷wld�y�ϲe���!S��i�S��t��:�ݨ�Lp* jx'�^��snSOJ�˯xȏ~��6O���V�D]����\>w����V*�� �(��ƌ��XfN�+�/OY���|
2�;��h^�ZT����᭽�_�*��AZ��6d��؎�/P{���s����C*v� #�4��LI\f2�?�+�B�+s��%;��g���_ߴ�u(ŲU�(�|�b;/7��:o(��!�o��&VA��U"�I�B�v1���d�tJ��v�P>��HR) &l^���'��c����e��>/0�ʅKT�@�P���&��5�\�g���M��N����Y>��M��F�]c	I�=�d�7Z
����oV�q^�sC�zI�hO���?G5'��-gg3|���Ԗ��7��<��b5��٠|�gp�n���)�C���SV�V�O��J�,�F4a���i�Qt�"dE8�7�y�����%����٬Y{*����:��2����W�ߓ/�{����Y4h��4�7 �-Jȶ��';�S
	-�GK�k{����E�3�i�&7�/�]��P)7��4lR ��J�,���餃��t_���f��Ǔ����� �4D�R�`��$�*�\�8�'�T.��IWu�Q���K��^��ms1�ɥ`-*�C��xks?�p���pkEIa����J��U��:��7�+Py�Ķ�U=�Ȳ%����L�-u~f���E���0�1������j(��e�!>����?TQ�����bn
������0����=;�����O����^����� �YǨ�U��ow*�vQ|.$_�)�vΞ(=q���2�z��T�0� f��Z�;椂{��$�;b8zۜU7u�]�[8W9S�\�,j�Un/,3��'�a�mY�O=��3����������"JK0 ӌ5;�^eG\F�	�Λa�_��6�6"����r��+��OVY��f��;��L��K�yc%�/�뎫AL�3���A���o�Z����_8l�5��ՁA�PF(Zx�I��o�\6G���Ɋ^�����hm!DyH����#-�t�Y�qc�8MyPt�*��f �#�櫌��|bb��/�zr�j��{e��T�,��{!�d�Y���?u���W�W`���E�3��:?��G�9�'�'ml���rꦽ �<�o`����O�}D����j��r�
� ܲJ>�j�~� J�Q̭��8꙰��/��5M��r�<U�쉞'Q#?� �F�� �Нl�bKzth�Ґ��
x�ð���{Lsm��$_�?Oh���ҭ�em�,��_q�f#���Qۙ^�g��z"���.�*$��4ämr"�_[0#��x��.��� ���|������C�-3Q����$r��/�Ո�e{ݻ�f�����ÁD��m������� Y��p* ǣ!#�.�i_J	�A��3+^�ĺ���J; CoR�w�\��~�mS�L�L< ¡���Z�0>Y������R/{���T��)P�Ku��v%-^�j���6�e�N(�y�;DسjQ�͚���X2��1M�mAK	
59�f6�F��G��T�ZnM��%B��Ι���Y�7 �b�N�x�a����r��d���Kp�k�fd\�*�����N���3��S�UN,�1��p72�I7�#�m����kߣ�@�1JHP��9G�єU�]s�h|�E%0�60x�*�t�&��D:G;��J}Q&�*ܜH�u�Ʊ�҆ԣjC�i�Dek1UG�yVd�$:8a)31�*]�ގW*p�Y�{��D>l��P�5�ĩ�D!�ґC)Wc@��a)��Uz��&��'��y���I��#1�R"4����$l��gV\�yElz�l0�MDS��8 fiXr!��xg?���45�P���a,��WJoMD����VD_Э;����}7��e[�l������D���)�4� ��4	��艨���.�m��r�A_�+M;5��!\�Y�mO��d��,��b#1�(`����@�E�ˈ�9F��>�g���G�L/�cRĈ�x'�,S���Hύ�_�Kj�1�cu)\M>L��D�[�<�F;y����g7P�Y��Q|�K���{n9K�vMC&į�Ӑ��i��b�_J��>t~_Ա A���ӂ�SM@4����aE�t����h@�sw��Ut'ٱ��PRZ*�D�ԓ�V���U����k�߾ϥ��������Ϸ���v5!�h@�T�va�f���n��{͛_/��/gf�����5<�gA����Er�·�A�rcH��^��Ƭ�H��-�T%�����B[m��Qv���>�Y)�$����2��iN�i�!1~���?��f�_�u#�����9L�-�����2��6�)}�>���}66��Ƌ��&��k�0�����*�k�|fdk� e�vyr���c.� H�9dt�E6��Y`�:WN��Gv�0��ַ\���=Y�o��6��>w�k���Ms��?�{>gsv�_���^�}fp6��r�.<���'�2���	���۠-X�9TL�ȠGP����fKǌ��Y٥�e�~?u`^�����Ţc6? ����R	9�H�^�IŜ�Z2��*�+��т6\+8�h��e(Q�_��at=(~�@Po�=�6ym���Ka�QR�ݧ�Ҏ�N�h�pH�E);�=?��i��EI�s�k�Է��|�o�H�g*C�_��΢F��y{c�궐����w8d���T�Zu��^gC}۞_���vqG-{?��ډ�csPw��T07ml>k��X4���KpH�j���fk'QU�ɷE��|�����ѓU��y�sw�� |i�D�X��{�u��o����dQ��pK�B�qF���E�^�=&�j��5�N[Y��^<����Ţ�&w���=������1�D�?J�i����2#���M0y�!t���?���?D����)UC8�(�Q�t�F|Qj ��e�~�P-YPZ8�Hx3O���L�Bi[%���Dͨ�p���f � �U6^��`l�Zgrѷ�{6_��B�W��l��x "�S�Y;��WE�yó�s�{�N=�C�S�
�V7f����o�ǹ���ZF��.7��wu?D�c"?�7,��-�@gף��i<�w9��-T�u��*��7���[Ȭ��rQz�ha�z��<0��]��"?�ż�oQLNwi����Qy{%rc�v?�RT�A#�����`�(+X��9Di�9\
u~^Bu�ˌ!��I�Z����f�DԴ
��m)�_A5烤�k�@�����r]�A�#&�I�b8��T�<L<i�Go�j�[D_Jsr�;�%LE��[���f�W��	TQ�KEL3�ni�Mh)�?���b�!	O��=�c��C(�����F ȟ(K\���g�I;��v72�^��ѪH/���Z�\0�u�ִv�$e��?��cB��@��l���Q�_aF��v�d0٘��[c��$d#����<(0w%��Z�w�_�X;_�N1���w�X��=��X�"Ï֛�g:��8 #�,��og� �7T��cHO��PF �Va8���R̝� X�!$�Zk,��M��g��h�l�P�ڗKne��)�M��{�ͩ�i������ٮ��r���iƦ�#�4�E�mb��s�xwE<0�楷�q�ϳ�#QLr���H~���{3���\�gmo�_3 �Fe�=#��2��z+p�)~�9$�]�
ӌ'i��m��P'-�Z*��n��y��%<o���^6V��0��>\ƸO�J3x^$2�vCO����<ԎX���T-�'���ߑ�5U<]�i�A�|�awڵ�5Ȓ�]V�٭Ա%8���cd��]m���Xw�.I4��r�}q.@j�ҜZ:�B�2O���q� ]�����������E%x�
�ߺ�o��}9�&��`E/L���I[�|��Om���7��X�����athZ���M���,ʚ�����ZV���sV�1��'�E���y�_�?���VO�R�B���sX/&'���S���>R	g�o_$.���?�9\�'���o�D�Bo��J����������sZ4v�1�}I����7&�g� �/,��\$s/�'�E�k��_&������5Ă3��b�S��JF!��+��4�桙�v�䘑��]�)�O��� [��KI��#U��3HS�(c_t�u8��m�&�)��:B,�2F�sK�)����'���K�V���\�D�,0�6z����Cvs7��*�?1䣁�[�C���-p���Ynəv�Y9̯ާ��

������c�T��d�|�L���J �K��j�����4��&�D"-���s��s^l�ښ|,a{ĸLH�0��l�:̥�0A��r;�Dr�5�֊[q�TlB�hw���I(�5y<��[hm;T��^G`Dq�����j?�_��$���۸�,ŊB� Z��6'G��<ڼ��v�:6Kz0�,� H�����"x7��KdV����v�<�A�
�aUkm��5�2��wޜr
+��6
��B�Yg��8�x1�&ǵ�9��Rsa%����Ԗ�/4_|��RL�]֔�+x�8�"n��4�u�r���'�LhT�uoq/�F�-�AY�0◀_�՜磑�wm9:�O	�Ͱ�{k����D�8{�=~\Ȉ��d*9�Gt�ߊ�)���b��|���9���.��L���r��$V|jQt����h�}R�A�B,�"ϟ���a�f$�
�ޥ �@q��0�0��g�b��o�Q�WW~�T!#o)�����W����=Uc��b;s5&�C'/�JE�/芙
���w0o}0���g�Me8���O�}f�����v�a���� ��^���]�>)�1��*����}���f~�J��i)�x������=��a�r`�� >���vv��1"vmk<�r���!�=��1#�ءY��[�_;^�5����(O߮tάYmp/����,���wf�R#��QAW���/��7ؤ��޸�KIO�ŉ�-_�p导n���� Oyc�'�v�{\�;?�,�9�\�n���ƭ��!�@��b���(9Ϋ�/ l"�4�(�*�=\_�G��8����@G��6֌���3��nq�)���,nv�ۧF��:Mvk�<9Tq�x�xd
��M�*�:1�h����k����Ыl���HiL]���Ŝ����k��9����H �>�	-w݊i���P��Շ�V����D~(�L9�俆o�}4� W��֍�5�'��d�y�U�/��n�(��Թ�����+���l�,�*�N���袗]�?�z�,3��W�$���j�Ym�'���[�*==R��{�x<�;��C�_���TW晉����`�
�M�[Y�ZQ����k>��_�Ķ�f=?��1��;m÷�{�l��A�#�*�cy��	Å/�[7�c�qQ��w�|mV��܊��s|=� 6��$��@�?�?�T��nd{�r��`fE��X`|��o컥��W�ͮ���67�!='C�[u�FFd���E�z�K�|�sB�3 ��<�G)C�	��0��7����wg%�c��P@�{�}NlZMIm g�N��L���ZI�P�)�u"���ASpz��"N�j���8����"qG`>A�}L��а;"�ׄ�|���^"8I)�)L�^��Tr��X��e�c����5Z���a��1��	[��:����CpZ�	g�h}2�������4��6*�>�X���i�is��o��PM �|g6Ũ,���;#��F����S�u���l<�oM)å�ىnk��J	��CۢC�ڹb@S�Ԙ�0�f�����BGx�&����X��g]����!f+oTE�*	�ǇY}������
m1f}�3><���
�"�]����h�|"�L� f���5�`�:�R���1�}ƫ"t	�]�r�9�4�EG��Mk��bH�Ҷ�Qvi��
�>+WpR�z ��4$�?�XD�K87��+��N�Q˒ǌQ+�LuфՊ��f͖G�>Z���䒺b;!Dh�.j��bdyU��q����(�Pߖ����4q]�'H�Kc�.V	�r� ㏍��_��R:�� �Rl3�X��p��Ic>�M���
���Ձ���]���/���:��w�0��,��#I�D��g�J�(�*v�n��),�ۋ����B'}"�[j߮��Q�Ұ*�z��=��R�ن�q�4}\���#C�����@;n@��GD�Z����]��X3��$� ����9ȅ�O��lң���1�u�m���`s��/�i��h�0�\"PV��J�n�X2B�P9�SrX[���G:���߇D8��^.mȧQ��@���K�Ǣ(!w-_J����t�T񂫘��y� 8�-����1�9�חs�u��Rx�o,������R�|E]X����J�?g�P�'&���	g��V<��z�?�֭�Q}���t�p{K�2��X^�x��a��i����=�|���������!^�g�aI�yL�p�������^�$�F$!�>o�Lva"<�|Q������i��]7,����"�j�7�?o�|��A|���^��\�����Q5G�d�ɝ�>�\��O��t6n�`�9A��[߲����OC���h�.wa��[����uH�#+�]Έ�ڑ�D�I�?ud$<��:�@I��)�9r�s�2��Fe8bU���	d�J	�2��!k���Z��l��'�bC�S�A���E<#�g�
Z�����Q<�#��)%@yu$�0���nK&����M�����\������3H�U���(ȣxw���gV*4����4ʵ���R�o�a��2�с�y��S�.݀��tH�+:Z�L��w�Q�~&���O��U��KJ�]g
�����L V����&@u@�݅�c��D��	�sbd����m�N�j�Q)� ��Bo���J�{=j����N�s8�����x��WesVC����o��{8��oݔ�x2�F�1U�LD����hƑ�%��r,�a��~9����	69���q��H�MwB����N�2��CY��p+�|�z)���T,�ɮ,��9Q�(`
�=��#������Bb�h�����c��쉱��<�݃a9��c�g�$�n[mL�Ǟ�sY����r�y��M\i�(BNsN
�ǎ]Vq&��	�쉛b�"+�tث��D��H��湼A�{����|����#�ht�S	�Ӱ�x,g�ꁚ�k��t�#uCMU�_V;�j�"�z%���=�.=�o$\^�n� ;�?Q�� �7y�z���@�]v�P�m�5�E�V�x/��{��c��G�sb�Q�x��7e����Y���f�j?OĆy�kފJ;A��Q}�;��|Ѕ ��GG'\��6<���i�����l,��b����X_��@��o�$��=��Q��Ȁ�A��ڌcΉ�\��:����[t0���3��/�4r
�R� M�ހǋ�El��Kv����8IZ�]�-� /*c�"=��73ꎪy�)L�t���);��zߖ�(���'��Jt���υ���^Nl����I��S��᫖p ����曬P��n�
�ה��G'K���}l1���~)a�}
��ӹ[���޺��M��Ϧ�C��������J$��~�@in����+��S"��zf�$SKF��K���l�{m��#O,*���?��CO%tJv��[K�T\�DU������RZ�%���((OE�_�{hd�b�p��$C����r(�V��T�V�

��?��0 k�*k-����^�l�WKUM�|���+}���jɨ)�YC,x�h�K�|�}z_�����
%ʋ�q�a����2���V�
�j�K$��|��o�n�D�B}r�F��+�;f��i5��S\r"Ue�g:�Ir�g�h�{����[}����_��Fp�4��{d\w�h��I�h=Ԋ>#���։�{�4��6�B���?eh.��9G0Y���Q��p=f������4�aeigV6�[�,^ԐsS �f\+�	)��6�HPv#��3�ڐ�B57�w��8�ӱ�ֳ� ��z���뇌����"���x��Ti�������S�*/L ���:\�,GtNI��_�H����g�3�t��3��ڤs��h��	�@�7��0ڏ����Y���Ek�G�1��S6�<�iIe$�Q����'������o6t� �[@�ҫ���ZR\��[�����q�eiS���zp	Z1�]�zu�'���������홳� ���C�Œp�jRb�c������~�j�=����ZI�PȾ	L�r��f]\�-�.R�#y?~�_E�q_+q��ʤi�'�ʳK�n����{�k�(#�5qNy��eq��T�f�"�
���O��u+VK���x����}`g0RY��[ �P3s��8�t�񏥱l���OHe���~�K�0�DFؔ3�#�毩�p(y���%�0�,����������O�u7=�k��$C�5xw��<��z$�jhA�k�ǅC��y̅�H��0lb-����!;�z
p�*NH�PI�c��ʹzU�O~�BM�Uv<^q�N��EYΨ"l�.7g4s�u��r����kS�:�6�Cc�;O�%�i*�d;i���8lЀ{�@�k�%qU4[*�<�Z�.��
�;ߊ�$�:Q��#�S�K�3� 6tl]� Tv�������'��_�'4���w9-ɼ�.j�ř:��1��؏;�iv�Z4K�m;�����h���5����U#���~����h�a+���ˬ�7⚇�)c��v��A�.���  ��0�߫���t����zh	p�ݢ�O��*#����<8���`��8RTn$��8k������1�a �<��`�n�����|�����S�b�%�WjILk��Qѯr�)}L����F�I�8��u�`7p,���� �@�H�mi��J�� ���s&��Ļ���f&WC��M��N~f�	@R�#thkg�V���$bcG���.3NoJ��}׼߫}�G�8���N��q�BnB����o�;^�{:�7�є:�7-|��a�A�B����z�o�\4lr���Ч�S�����c]��㥅����C��U־��|+6@B*���=Y���l2MA5��a����^b�C��M���8�3xI�Ҍ��i�~z�4PxM̭Zݺ�6lO�mV�&���O�V�R�+�(�����Ψi����?"�k@Ե�"��<d�rB�B���!3�z�Hɳ�v����13
��kH�{lW@Yz7��SX� ���s�3Ch΅vm��n�n�R�?��˼IA��r,u��g7,����E-8Fgz�dj M�&~6�O��%�^4��G��L�\}�)�����ɔ�x~�O�$�X	�M��	W����
�W{����Wv���` [�䋽�([���n��X~h���F&0۠���	!�~~�d∯���xtg�bB�O�#�������Ҝm�����o�0�{9=�[Q&��Y:<�H��m0zխ��WC%5[�r4�R��*!��> ��uv�v�k��Gf˞$t!�<h;���	�f�q2ƕ*��G�hN̢�M��\lh����i��V��B�%��Ϩb�s�4�1Oss}�����@�L�SF�����(9�˖�:ӈ�6nN-tL>�c^�R�ξ�I���U?g�r�� l���<"~A��F�����ˁ��w�����O�z
��P����	�_��z�f�>���Ǽ+FA� ���og���&�~*ÓE˹b|'��o�����䎾_#�+�Y��<23a���d���LM�gC�%��`r��y���6	�&q�Q�S����jVЊٙ@rRf����>�&�:O7Հ0t�$�Q��<�^S-�K��N|ˆ9)�@���]�5���RP<���|��M�J��O��%|!���zɾ�U�h�0E�1-J�G0��5�tF��+?/��Ak����n�S�*�i��x5�*n��ZU�v42q��������x ;�@��v�Z�O��Op�M�H����,
0��Գ���@,;Q܆.MN��N��'o�e;p6>�|?چ�/��O�C�N3�l�k�܊��f\|�_����3�q%R�5�$�����[�I���ǰ�#������=�2���[Q5�<^j����<4?��UKU�N����Z�dD���=�Hb��70.�[E^�M�f:$�h��
�+�e}
�D^.��,~��`=��i6:� �Fʍ�F��20��炗��Cl	��A��6�� 81Ӓ�D�?�ٹ�E��g5��2��g�|�	jc8Xy̐%�-#	�a�����|ؾ���b�h�u�4��[�ѝ����Wօ|:��<��7�G��BM��4��o��I�B�-Nm���9���8�s�� � �I�L�Жz	�6n���hqK���70`��n��M��1��)*��6���^�D�C[�q��1�4���}�CԚ�$4�I����F��`�2��"۪{��|�u"`������~`�s�6�[�Ư�1��
��5VC[�#�FJ���p#U���|����r����m �/=s,]��+bY�0Mjw�T���'l���ha	t6�RW`���*��bb�eK�7���pA>VD����x���h�w������[��r�������j8E���;�� �fI��Ɵ��~{>�I�o=ԋ������]!��g~�/84]QÄ��4��7=|ྲྀ`�q�q��x"'�p)����D,R�tT��R���TNz��d�/�����g}��a�W������%^�*2�-��^!sj�ĉ�x5���s밍T��������|��A� fk_�~Ļ�\QA�8��ާf�9��N�3-�ɶ�����D2Wtu�q���)J	~�!E�F�y���7Z����|eI�k���Х�ɠ��W��0��=�g���<����ȿ�4�Y�VSN�%)��m�/�M�M�E�Tԇ�kgL��%�>\���.�KZ��SU��ֆ�2N�m���"#��w�Uϊ 8��j��r@a���7��ݵ�}�0��A�r_�Q����r��yM]�4��Q�ж�1�e��LVy,�(��㍛t[�1�_u���R<U�։5 �];��Qu/�=1E^5@�" et%I@��}1m��/J`���K�j�!�
s1Zσ>Jɝe�����>��L焠���<�G�MH�#��c������:����U(y'E(w�2���1Z�3V+8�v�~�i؉�f0�C 6�LN�'	��6�\�g�FF�M�	���i_�lMݺ؋�O��1�bKW��E�"���)Q��rGg�R����頉;�Pms�3�L�&!�_�a�~�v-�@4U��J���������dLuۂ�T{ކ0��d���*�����k�U+Ol�)e$s��0��ɝ^���.)	��{m��?���K���S�r�w)�n�/�+!1\��A[E��.��b5*���ڴq�`���()�Rݙ�x*fP�Ľ<�7�0A6�n�u1�M��(����g�]��2��J��������7�
��/B�����n��`(��e�J�
@��<~�&l�(�R����P�4�������w�����|K�#'�t�o��-2%�jH�q��M}	�R]��l�x"{[3u���&���1��:�[@ͅ�E0"m�_�	G�߬C�L�zޠ>�u�A���I���Elݿ�:w��m�*:J��h�N�tPR��V�Y�m ��Ѹ=>k7(�AW]B�zV�-�t��S�\��G�a&"$]W���&�$Տ��i��)Ԙ{��d�	��1��
��u� ���n�6�PQ�7ʬ-v3 ��r�V���2<�6n2Q�p�����պ�l`�B���4I�����N�Ԝ48�13ߚ��q,A��B�����$'ױG.G��E@��0zץ0/k��q�,�h���f��m�H��=m0�䵃�XV���z֕ͪ�d��xn�
�"y?���b�*m���6ho��������rZT�	}�yD��}�^�8s 	� �UV9�)*$βA�I�l,��]���O�ɿc���N�X��	3f�G909C�`����{��H��;,z	?,	�8=x_���"��gG�(}x�q���Ȱ0�;F�/�%	/|�p����P���!����.o��m�
�X$~�}5Ñ��f��3֞d�N����*Uy/2�Vm� og�$}�vn�uH��)]W<�ܻv�o�2��7B�#�&y����������ю�eg�3w1�c/"���=1�F�v���9���K3B����ҹ6u�� �%�l���Iq�+��v��KV󾣥�N�Z�����1�`=�h}�'�IN��aZ��ח�ϋ�:�����R���d�8���O#n 3lUaJ�>�)�P�z�c�^�B�OFO��ɹ��]	���B�n/�0����Rk��u�62��t���_V��t��q�W_GJyr���}�V�.[�#��u�����K��&���#����|��e�����~Is� �������Gˡ�{������3�Cy����O����n�m=㦗d����.tJ����+�H�/1!@���$��譻�P�����T����t:~Lj� ��q�e��Hw��������s]$ϒi��Q�� ��̘����AqP*��W���P�&�f?������F�%�>��q�3�s�c�.#���̮��7~���U� 5$�k����T��1ԚPt T�R-��Q�7Rs��Ӟ�޼�1��uz�:겱^���P0�
+��ƭڅ,!�,̷��K!`�u�����0�ŉ�V��+�8��b6���8+jz�6�+@|;����5��=����jG���a��cp������Ԋi�?-�t�ڢ�_��D!�`�O�i[���U���Q���%P��(���Є~�h��j��!�G�1�;�a���[���op��G36�KK|���J ��t�ÞdE{}@v8���g���见)ƾI�b�S߯��k�V��L�TR
E(T)�g��OH�j$J�H"�V V��O���Y�[��~;�~��ƣ�l �Q*�1D�~��G�&e/�P���z)�3�q�_&�*�>�V�����9k��� ��@��%�i(iw��<��w9�)�Jd�̱۠�U\_w�Ѫr?
��׏��uSi4�05���	��Z��a����:w�w�	L�֭��j�ˮ��$�L��vw��4��_�\��M��RO��S�cP�$ă�~��ళ(��2z+\��]#_��J���V�����-��BY�����z�w��_�x=�Ƣ��3�1���̴�����\3�|�Z�g�n��B�V�ө��d�!A;�7������c�.�qO�z4�<- J�b�4��`����T���_:�д�o���>�f���uo򣾐gd"@��WZ0��c0xU��HҰG�����1����GFeL5��;]/8 'bOQ�,b뾟�T��y���Ic��?�J[�٫Gǵ��B�����t{��S��ܡ�3C�;�y�W�H��8KsW3����lT,;(��0`T���{��K>-�k:�b�Х�E�LkL�V��1�)�W�x6eqRu���!�h�b.�4���@>�_F�R,��M����~Le�0�J��Ef���Zv<z{���o�Nc�"������P��ƅ�Oзb�/���`ζ�+����9߿V��mGzh��z�?s\/�c�-�
~�E�73-��FA���A��p5!�4��LI�҃����.��(��W]!FY��^�o�R̩�rW��l�������6��B�q��0��������f����A568���a���l
J@ϴ��6�ZU��]X�;ɤ�l�ٸ_c�>t4�[�b�Y�w��y�X6])��7J��X�r#��X��mɺ4��&�M�EhE�+e���{�����m�l��ӭ�����o���pt��aַo�cM�:g��ے���!ʵ��OE̻P:��r�m�ǻ8�As�+ $�K�/<�"�6��!���W]%��r�J
&��{�$���z�~�}���=Y��d[��A^��Q)w��'*Wʃns�iٻ����^�WIa��y=%<��Ow;��f�3qRJ�n�pټsG �\�
U& ����r�%5,��W8������OG�[�4f����H��.Q��z��)��~~�
-�1����
JU6l�ɿ�a��b���h�/�]�	(6`�0F��<8yS@��W��_T�����C������9���04� �?���QN�~����/6���NՄY��I�lE�� �P��O0��-y�,���ՋL�6��`�1)�*�Ќ>˽��D�C��G�ñ��Vl6�
��sz��+@2s�ʗ���v ���{X.�
����3�:��>��/��W�6�51u@N�Fc��u7�DtA$���LP�bL��v� 	a�fs�kyPS�,��ß�>��]���n�'�bK�Gz��IG%��ہ���P]��V����59ؖ�;�.�j��䃛�?���jo�����X>ƈAa2�q�x�RX}���23bIE}N$y��w�R�QcҖh􃁋��2�*��Y��BM<�x�ط�"&&6�$��z�zeI�}�jK)v���wm��u����o�F
l�Z��-,(X?#?�rwr��T�]�{6����/J�~a^�/AmN�����]�"�ItMޔ�EQJ�>�j�knӺ���M�͉�R���N��ll��)J{x����A�?d-!G'RA/4��ڴJ��&�}]:3�b����˽a�ύ��f
m�SO6�k�Q�\@dWf�(
���J���kPtņ��4r{��ɯ���.��i~�_�<�� }x����,@����|��Hg�˃9����L��5����F_��k-/ڮ��Uͫy�R�ȥ�oc�W'o�A���謪H�����hz���L�C�	�/}ч�%���F"����룤z��*�`�u���ƿ�1u��k�4���ʇ��
h�x�?�v ��(^��k�D���IQ\�Vӵ�!����Hp�K&�������h�k�b�Ƈ�n�~���TS7,�ж���߬	I;a�dx��Z%���\��)��v�7�v�͸y����;wݢ��=�D�ډ#]Ln��zn<��i�/�#̷�þ���o�#����ۍ�?|W^�W�p������t� &��zJ:*�</y]-�{�/J�e���+���N���|u����5���C{���V5jUa2�y�t<ĵ.�%��T��1a�8����?�]�YL�Q��t�b��I���|d����0�!�9w@}Nk��9�媮�`�G�����?;l��39�v�wN�L�T�����T�ĸ��15ueE�W���\������f�RM;b&�̯Pk �ס,�5J�̌�ޒ������ɚ��Q K���~h�K���3���O�ҩ�R$N1��L��b^�<��i���9T9���6�!&�
��p���2�L\��L�]�t3Hn��⨩s_ ���/?s��q�{��MC�܃��4AI��Ұ�F���.-�J���XnE�k:�jժ����|��FⵏAm������Z�O�;Bpf��W	����U�����҃�{8w�O�ڋ:R�a_ /��<�p$��C�l05�[.uB?���M�� b8.�_\b?����=�l�4��9̾�Y'�.�N�bk��+z���2���ʙ;�j�2����"�E����7}�����ԏ$�ٞ�gi�/5�rO#�%q��4?lX8��J{|VҌ�\�;�P���7Pw�*CYH�����elbti���>曔?l~�D'Q/�6��*;���َW����Z�����+��%�H�d�����>��ī�`�Zh�D0���K�*k&�P^NQ�W�ȕr8��.��<��b���z-�P������xj��~
-�"?�A�=�҆�.XꝲH��뗶,\)�t���@=�!�"��c�Z�Y�z�nӄ7��]��g|0����'<׌�=�Lu�׃��A�=�6z�oH49]���ޮ�;�L��@��r����Î����4ڔ�����Jk����^[�x����s��m�V	��WTK�[E�dQ�3o���	�V;���^����<F[QφN���c%�y� ��]f��ii�[�M���*#ë�t�O4�'�h��Bɞ�jTY���";�s�F~_Z:�ܦ�;�k>��
�Ü��!��w�i��ZR?vE����L���	�����o+K�")�x� �r����황��Igb���ӛi�BP�~�A��?���{&��{3���0�x��YgO�sEzѺ�ӊJ��t��̾pRmڦ2�QD��T6T�j������8�$�D�����d>.�b���G��6!�,-�\��-��4�Ya[q��^�ي�,�B Mv�9pͨ��b*n���$����M$���|v�>-��,R���}�[���yh�g$1M~��ٌ��:��)�8��-�
,�.ĸ�m���^��&p���M%3u�o"��F��=[I�!�$��٘(�P2�L`m�O[��c{���ء�Y�Uk�G@*?��|�^�@	��n�U����ɡ��3qx�>+I�O����}{zOZb��f�>1}����1�5���@U���)RȣǷg�\�y8RD�M��[!5թ�����Z;��;;P��y�J����`'q�aM���',A?�����Df":�.�lQ�X���@Nc߀^,�,يL�h*�7��ThC$ᣐ	����E���u"Y	�rZ�6�c��N\� �xPK1���|N�n����͒�^�cG�X=�����ƘD��U@���H쫦��A���շ�5�a<��̕S�i��}岤y����Ks��X8b��:��|��c��@j�	����G�1�4�8���$P\̄�QX�Z��8��n����"� ���U����מ�ik���4�%��}/JVc 	5��8v>Y�&���QE�ilN�n�8J\Z�^Ӗ�(F�[\�3(+��7���UJ�ϔH�0�t|�Q�W�KOF,`��n�4z�{,@�Wz.lG�6���J��&��I5q3Ed�$=�7�ze��K�����a |9�v/�tpvn����T�ʳ��D.��K$��o���{������M�2uT�Nz}YlD�L�6�AjyC�����������m����ھ�&)����F�iXd�������+n��Y9v���xV����|���������"��
Y<���%��|�Ĉ��eHf�@��u�c��N��ż�;�_�M4�D�]��\���m��pmB�Pw<�� ����3��^\D��/<�;-�2	:����3�+ͳR�ʜ����ɂ�^����O�h >@߄�a����0"��v�E���KJ�ӱo�P����~����rPXo�7�R�+�zR@"����;(�KhI�e�k6~�JĹ.�%m��t]MXb�@�_rF1�X�l	���t ��*~��0B줐4w� ����<A��Ҹ��nKY��&�p�>��^����1���>���6'o4<���
`4�ؐU���]��ܴ@{�Z[�F��R��\�#G�a�����;OM�ۅ����w<Y��h��&37Q��U���|C��6�/�G�M��mF�u�*�O"n�N���P�X&��vr�ާ|���Jq�k���-�r֗?,�փ!-Tm'�rM��s��籗�Ӭ%�*PݕԖ�Q�l�A�*�F�![�k��(�	hs�AN֗k̠�"�:罍�1���穧l��V�k��oPJ�մ�^D�o��<'B�h5M
.ۜ�5����%-�����2gX�q�j�c������@:.{�l�o���)/��P󗄈*�s��t�D�x��)���
4�}�tc� �9�����iim�Ig\�|iW2Ŀ�h"���ޘ��'g.~Y��X���{�C�Z�]��&��t��ܭ�`��H^�+�e�d��m���vڬ�%�%�Kx�@R8��^��jZ� �s�Rw��w|��:��-�Q�D�ւhN�)Rv��tFʄ�,�@���-��3��oB��=�a�m��C_�g���������.����vq�ţt�#��g����5���E>KK�ttkds��*MU�.A]����ˍ`�i��^�}�	m��/�#b��z�4Y��TØC���L ��3ڇ���Ty@qj�hu���D�'+jߠ����=A�y�&؆�24���?h8S��r��t�{pɱ�̓5�-���2�} r+l4�*)m�ׂc&�*�ŕ�9~�99������ՆNOŏ�;��a�;.���Km�%h��2,�+�_��I�6���+!c_������3�A��QU�>Vj���}V���� �<e���{%����mj�������&vV0�no4�	Ͽ�e�i(�A/sm�i�����eEqD �"2kŝ8��[�Ϫ�9�Ⱥh��d�L�hQI\R>T�vt�G�2���
����G�i��RB�3����!w��l(�a��>�h_���~�>��ޞp�>��DH�O��<�fl�6��8<q�'��a+�b�v6�B�RKoP|�PO����T$5�����z{!�|1"94��"T`��*f�#�t���_�W1m|�ݭ(�S�CM�}o�p��(v�����:��y�1-V�*c}2f����,=����Oy������k�ȓ�*m]�JJdH۱_�>�$FmpVbE"����y�E4�7��e:�&g<��d�={��U�����8��	vƣ���C�
�[��쁥_%sG>v�
��� J�5��T'�=*7����|4�g�b�̕����Q��uY8&6����ig% Q#�~%�E��GW���j�~�V�}W�9??�����`M�ot�*�y�ڭ�셫��&��@7��^/��N45�����
��R��m�yu����p�	��_����@���2��3�i�v>29��Ee�l�Ys�@u��G��3�Xt��Fq��&�7��GT�L�B�x����63�ޙ{)�v��V~���Ss�D|+��`��k �.m�{2���^р X���E�"Z#��,�ϗ\��n���`e-�_���2O���C`�Y72sT��"�Mݜ�&]L�鳑q���BMW�8�/�ϡ��x���쯞�6�N��'��ę���Q=K���+�/�G����|���r#���=��Uk���3d'�a��v~]o��8B����J+5�Up�f! �Ӛ'"[w�u��J�sD��F=p��1C%��,���� �"��`��Q/����c��9z�m���r�Ӈ6I�	��U1��xbLb���G����4��Kw�V���]� ��]Ȭ������[���q��XU��a����]VpIz���x-����ڙ
VH�_ÏA˦K/�]�!�{T�� O^vۗ�{>5|���r�Jg�M���7f�Gǒ?���2�[��z��4~t�+�h�툫�J}a�#��0�(��.�_��WQ��O������?���9��>�Ќ��a��?��B��s����╋Lqr���sB�۶�s�؎���u��r)��N��3��9���_�V�<WA_Z,����4��.$Pci���M�����fmF�:+^�uG;�E)�ʰ�"]I���=Vr�QH#ީ�aL���.j�/hAK�&q�9�+`��gcx;�E���\k-'�$�S�B`��+*q�ح��&���+�b���`z<�2r�*��?��w��'�����d�ǆg{��}���C�V�tv��K.ѥ��^�,1��5�@P�`#�rv��.�et����MX�8�0��%�0��Y��1>�Q����%l�L��Y�F�\@�����y��D���`vC���f��,�<&�E���M��?�G���e�w�s�0X���K;z�1��-	�>a�M..Ӷw �F�^����#l+��>�?}\O]2�%R�����K���`�����4r�S��~C�	H�5��ɗ�	`خ��Qq�V?H�(��9Ό���8��~(:�]����$�_�P��ˑ�A���h��(>�q��&��=cy��ix@�5���vEY��~������U�!�ܣ�J���aB� %�M�?�qA��̖�X���^rb��z뛈��U�82(j�w���po���1D��F�xxk�r@��}�p����O�0�X�%#���{��Gt����4Qܓ�_��)�b�R��1
�!n;ӆ���l�C�L��Id�u�-����k�x��F~F8g���@<P8��3h&�+�ev�[KQ��5�s<�-���S��(������'��\94�:�(����3&�]Z%Te��!9�cח)>������/~��)��a6��5�*�1묌��[��w7�س8(@�Bu5��x�+�ǀ$��l=�w=A�r�) d.��QC��­n�Bx )3���� � ��Bt��U�����H�@$4&�ڕ��
�NQ 0{�c�X��+g���N�i��ns�ȨF�\���"�h�[�F�&*=Y���Nd1'���j�+X4��!���<l4NL���汿-Vw;j�pJKܜ���bsdG�t�ɗeѱS��;Q�A$�鷬��XY����5��c��6��Bj7x��B���)#չ�%�-��╤`@P�!�LG.�7@���LQ�q�I���j�r�3�(Q����zJX���2�&P�t��൵]�� ��n7y"N;v��;�'��D䈪��J9S��@W�#�	�A'NkV���w���^L�i�t�G�~��g��b�A	�^�������#�	V4�/�^�e�}RBʑ�/�0+~�R�Ot��9.?�I.���| �XƂ��r��	rx3\�FY��8 �{s��`��`䣁-p�f��;̹h��O6��*>��Ǝ�}g��~Ϗ{����lpzK��$�[mM��}n�\f\=;Q$�`HU�'˓ZKBMƾ?��'r �A]�~��M���@�ϣ9�Ɠ��j[^���_Z���i�q)ۈ�ۯ ݎ��^��S�v��g�&ޯ F1���S���'�=]<��3y\Gݹ���D"+dՀ+ThIn�nb�ˬD�D�*�j9�`�Y'L���Z���T'�����ߤ�E� ��.� `!l�zұ��@�F���i�Y7@f��Ȧ\DH�h�j������g	�#�r�"f�0e�˖V��;�\�����>��\cg��,�t��	*��I�XF�ޠ�5Z�J��g=�R����Y�<~�E���>V�ץNZ��t� ��y��Z���_�VFO�)�n���Z(��iK�x��F����5������xC�\��6:d{N�׆O��q���L^Rr���+)U�r&��΂�[�m��������/i� u"]��!ZGr��M}�6���ڛ�V��u���|���0�6�[,Pۨ{}���֢{K�ݞ0+V�#G����D06-�)/���2����r;M"��_u���S���8�m����]|
دϸ�7��- ����#�J�'��%x����y����K8rY�}?G��t/�}k��؛��VK�'���Zhz���v���������v��}��v�+{Ql�G$��k{n�Ņf��cGP7'�R#M����r��p"j�! �d���������h���r`�T@�VPT��$�\��l��sB��͞����P?�𯙫PZxޏ	 �wOI�f˴Z��*�i֒���0Op�X>N�Y�\4P.��};v?-����y �����F<e�͌�k��I�$;����;r�7���5�R�ڛt�g*X���̰8�W�p�)�
D�%�^���?[��l��y��$HT.���Q�mFVV&�~�!(�y�Ĩx?m�͕y|�&���qa�)yf/�q�/O�=q�|)A� 䁰�G���,}a�9N\�}	�%�KJ��a/��l�#��r� ����P:j}�3��D�ƒ~�ۇR���Q�-�\Â��HE���NM1�!�Y�G�"춽7!k}�0�%@�xQC犁J�(�6ȕ�^]L�j� M����=�&#-ܡFl�c��D��'(�ht�J��["���k�J��[�Fa�
JwiC�{#Z���J�U`JCc�3�F�\jP̃y����D}k
j����a{l��?%ש�Y6"�}���G�E�A��Sk���LV�>p�`Xi�����x���%Mw~��E/�r�C}gG�=����He8�O�������`GFO7]B]��3��b�MZ_@��:u��ONt��$�u∋+�{E�9���gei]'(:|
�*Cj�Jp6���.>�08X�|.��<��4N�>!�~��vu��QO��
��̫�21�#+�Te���M,O��QWfRz�~A�RV��ğ._�˅.%��LVgXh�XM����Z�^����D��wL��@	az��33����VyXv��j�r�	vy\���gz�YD�+#������
8��]x���47H_ B*>*�N5�5�.=���]�tڧ6�Ӌ�U����j0�] �&m�Vv������I���^Kjp�E�u<���N�~ �H�&�']�f����o��J:����	A5�q�Y�G�\�����>��jki�i�_��9$�cw�#l9�Y�4��1Ǟp�cZOksn\�1#VT|?��v��Q��Q�x5ީ�C뉥)<�hђ����� h	k{:�s���߃��j�(�s/4c�	m�(�B3Js��Ҝ߬�.M�FD\���,��������FB��J ��ێ�,��ٱV֕'�p���g�fhD�i<�����r9�E4
��Nf���s P:o�:�$PT����|V��!���ind� �Ɉ@.���
��D�ҺV
�7?5���y,5T�*V�_9g���miҊ.w���s�<E�.���2� ��7Y��-v<wi�r��P��|?-����ĕQ c���]����b "���]~�o�s������e��뇊`����_�4�cΟXQ|e�P���nEډ< �ɲ�o`Z�:�I���`!�ŤC��L�FA[<�U���ʌ�y�Z��#��!6U���	�[�	��T����eU�rl� ���FX����b߸� 0�q�(�- &~��L�t�˼7��}e�]�aWZ_p夎��F�	��Y���:es�g�����
.�%F
��c��A4��x�23��֒��_�]�uu�r��8�i�aY��J�M�C�	t���f~��q��m�Z�	ӽ9ɼt�ܦL�5	8��1��^f�,UA�f�"bpb�f}o~aVC�u{��������&�v|T�k�8y�F:*8�
C����"p�N��ۙG�eELT}�冨��Ǯ/-H���
����ͻ��غ6뾊�����,��ͯIIhz��>��ǆ���h�x
���	>)to�d��g�B{��jY�,�*'�y��~�'uŢ#d5ݸ�S���.��/�v��O=o�*��*��x��/����T*�����L����A���ޒ���+�B�'���V���֔M��<��������
`�"��-��^����`��|�ݡf�`9�0�Z�{P�M��xC�.ʘ���6�,�)Q��R����;-۹j�� �F��d\�$�H�uJ�%U�\��\����R�����8��N�(�Y�v�fV��#��3���8��cj�W�@-��b]ד�t�N��\�H�R-Hq�j��3xÉ�V]����{�p�H���!Fu0d�7��p+�vB��S��O�z���0�7�q@�LZ�O3��6�L(�`�����C�bN���������"2��֨��%*5I ���F{�0�[�t#�i��pԢ��X���d�=qFDy%R���֨�h�M3XR$�_L6�M�[�]k�B�{�� ;�,�ʬ���<^l�n���_,)��˞C����W�$�8�=FB�o/>�I|.��I���k��F���������@���eL��L���У��G�Է�#:�)�P񈜍*E$x��<\�����ςy*���b� x>�ޤ/{`���� ͪm�/!����4�֗�/ni��N�x�l��$����ʠ,�P�3V��x��z��p{Z��u��E��HZ��f+�Ɲ���dw:��ԗL�1�|��o��2�Ϛ���-at�� ���6���E�G�?����ϊ����@��I_;���"\��K��a�,���SWH�fuw��9�f8JVۉR��G��Qz:��V���EY9v�e�H2��&��a�9��
�FGBtEJy�����n������:�g}�����z%O+�O����i:��}pt')���wG��KT�r�����ul: E��������Qz��N��h���a��^�b�h���#0+!�g�4{`:Ե�O����(sV�t+�� L�7�G�X����_���$H��ci+S�g�<i��C���$elA�w�����@}#�-0	���B�d���~�pD2��`+Z3��vX�k��T�K��ط�V݃�]U�cGY����5Ģ�G�>S�h����k�`��5V<���m+1��M�(����GιTi_49��D�ҥ�v�$J�&O:��ւ}�ϡ����1-�Y�����X�!�y[hN߂(��g ���0��sQ���n�ShQQ���wT�yÞ��x,�MT�Քa04���̽�ҏ;��5��^�� �U�rӬ�}�Ftsb`�譢o��KW��a�������.�VQ����I���ۇ�F,$z�a�o�Xip�AdO:NP[�}�k�τ&_�dV9����h�.J\��N��gύ�ݹ�I ��ی��m�E��p�tiz�u\�Y蔹�=DA�%K��y��WT�{��D�7κ��q� ^8<r�x37p�����h;wS�:|���>8��5�v%�2�.�Q)��`V�${��Vv��AӁ-��a��%��,��tԟ�'�	���:������/�Bxo]���ZR-e��� z�IW�eTV��O'C�1f��Iy
-��QK
׌��{_2��^tZ��b18�Cg�� �ě^��#�3�����/�l��2���pl�bb�_ ]�Ǽ3��U3����o*�d	;U�@O��(��T���4}���MϢg#l��8����ث��OПѾ��$FU�^F����@k(�[��r�U�_�;q_����XH����>l��E|_:�@3x"=�+����X���f�\̹=.D���p)�'�Gs5����Qde>��ܭe�otﻉwi�4�Շ�ro�P�,���!_�	X�������͔���U`���_��P�}�� Wk���=���cb ���0��P�t8����,v�e������w�d���;�ɗ`m9`��DW����[�x�H�֘�?�=�gL��AnD,&Yx�Y~L\�Z���3Z"�^f��OH�z{��1�b�'q:����2'�x�K��M��ى��QӖ�TQj��t������0�4���2!��\bG�.1�Oa��O����i��W|a��n��15�:n1�9�-X�*�mY�l!��?ըe5�0 ���/`Y$T�D�L�-��+L}�7�t�_S�aN<{�Q˚�e��9V��>4��j'?<�Ñ'<[G��Y��<�D�}�檊�2\*պىq5~'�e�E�����*x74PXe�etըZ�5��l�C�!�ũ�ci�-䑬z�B9�R�U�Q�@����˾�!2�|b�g��	�b�dԣ���
*�O/%�n���C����oTS���+�%[i����,215�}߬���d8pe�d����$Y���K�z�$�F�Q>*Zm����s�:]��aD�b��?�@u�'&��.���$��+B���_2gИf23`}GY�O��z���G|��Z8��K��>7#n��U`Y��0w^�s�̵	�!���WcT�UѼ�c��&���?�MIs�T4�����
mHrޢ�=�0��O�>.�͉�� �:�=YO��|�o���L��3Q0v2C��ό�Eܾ�l:��u����eo�ex����g}�?�*7Yc��Su���J�E1�{��:>J-���'�_j�����)�y�lSk���e9;�T,KЦ��Ua��p{=���Cլ�]�3-��)�֑P�>�m��$�82�d�J.km�h�Ԧ{) �B �Ų���.�]�{so�����_�0��%�ؽLP	�� V�`�%:�u�C�ܘNa������Cg�I�������;�JIK��{E��HK��c��@�<g��q��P^E�b�c%w���Ɗ7��]��W�T���l�Sw��>^A�r����B~�p�tH'��WW��\�ob��1����j���MY�pek7���,��%��g�۱ g�B5�&zާJ45/|A�P �]���l�'�ߨQ��O`��b;f�7�\���u ��_>p���4䐵U�{��m�/Q�g��%�9�r'��E ��ws^�{S0���V�k�y�����RbU��j�c���82/�5�R�è�~��u��U9����w�6�<�u0l��B�u�{<M6Ul'4;�ì����C�{��<&�(ЧsI���V���e�O�]��p���P-�� �ߝqbM��a��7[��z~|<_ϼ�Z~ƚOz�-G+lj�U�9�dm���5�ax�_|��������j��N'{��E{�}QyI��3������h�sv��^�e\��e}S�:������N�ow��@�,�Zb���{a(d)"i�{��r�}��O@������[0�Qt�w�����*o�&�gE�	��L��v�n1��s�Y�Z��b���>��Ƕ�r���ʃ5,���1�4#�ʞ���b[a�����^ + ���X��	������L�0h�d_�o%���jL���sA=�~����y9���Q��Lƾ�#Z܌Y�0)�&EP����OE9���(qϔ��c��0�)�G�X�m�2yO��q��W����%�@���8;����!%�,\��F�Sm��.=�3��xʧG#��RZ�ꊕF������~�|]�4!���h��A��϶-'�p����}Ӝ�������׎�NC^c1`x��K���H������xդ'������[���6s=���lМ
h��K�H�Yc�u�s�}�cS���Y=~�s:�;H w|G��7�Y��U��m̆?B���T�K���J��Im��z��sQG�O8D|xFU;w �bu�N��(�&�NZZ����s���ӕ��?�)��ç�S�	�D���d��i<�mI�پA�(kt���nX����TdK��n "���Fby;�_��wJ&�����ط}�cX4,q!ڴ�*���q�T
W�Ȗ�-2�)�O�z��E����<s� ������*���HD�2�';�-��%*+�m-%{>�H���*yv���4�L�G�۫(%m��rBQG���+��=�`�<]�*@�w�0E:ӗZi��z�E�!�OQ؞z{�֖dZaS(�������M�\�;��X���Z��(Z'O�j�8����c,�����x�ٴ�wᢾ?%"��(��6�hY���� ��U�`pF��8�eX�%C�j�
��:h�(�<pf�i����Y�؎=�3:_����DlUw�Y'��m[�1�����/;��V������P�Q��rpF�[C�BsO�K�༻̰���{�';.{]�q��G�tCV���b���: �2����ڨ^��o�c�׋v`T��ÿ��x����սI����R% r]�����37��߰5G��}�W��ժ�P�n��R4�$����Y��	�NK��q,���F0}H������͘�!�Qo$LՅq�����a�����?�Z*�:���S�v
dJ���Qk���GS:�=��١0�U?F�8�z��bb��,q&���_ MX�!�ˍ�݄�v������?�;�j%! {z~"���7��j����+�{��?���+e�G0��;6���	�%,��ԇԢ�bSI;3KnYК[�/95�$�%�5���`�.w_x)�'�<�o)�j�pP�!{��v���wl�����նN�>�#��1����Q"��;Ӳ�X�ǋ?0����A-#E��G4)��c��B������-��'o<�}/�<A����`RB��h~;N���Mͷ�ҥs��+���o���\�0�m6(����O�R��5��$��Ǚݥ�](�Ǣ1��ǻ��'�6qth�#y�i`�GGd�E`��9m;^8�M�nP�����3�K����|l�yZSc��鍜o�<p\�n��_�*�t	�$���u�$�&���{&��n�Ң�E F(�)$�	V�& *�^��'+�q��r�S���=+�	��>>���m�����R���_GKm4U�S|�.$�V��"��?�/e����|�g��$~�X�,w�9���U��	���Z�CG)��P�-{��݇5��\��B��%�^0'�g]Ǔ�x�$��s�L����80����"/L+�1H~���R@"�JŢ�<�K�(ֹ�<Aq9�����#�!��(��5��͗��H�,���9�E�a�Q�W��J��#�tA��V<I�#�Sa�*��F�%|�>��P��)1<����j�+״����GM�v�0���D_e���È1ݸ���o�0��������X�3f�z��l`-��9L�3��N���G�b"�Q�̥m ���� ���U3 |:�]�ګ���V;���a�0����1���V=X�+��?�}�W��&l�$"F��|�SK���&*���Hdc��{+��)a�dX�-F�~8Y�T %��s�pɥ��1�Q+s��Vx�^ l���Z���a�����ܤ��
�Ȝi�il�#x ��
GЀ73�� ��<1�������x����D�g��*�tL(^�yH�<���Ґis�o?Ƨi�'�Ȣ��[tm����?4�C��eI\��x.<�ҫ��� ����-^R�Z*F]RS1Zsb���,���s(8�$G)[$�C���G��5�t���V� ��^���H`I�eG��?E6 7ĕg#���68=�Q��CA/"N�j;�U��C�Y �|���'^<�3�+2��՝1S���k�NE���D���7e�t��3�#wE�m�5�_�~A���8�	6G���`-���7~3��6���Z0<ԥ/q/��5c�Z�?B�^l��n?��>�p���}K�X �d,R�(&zD�	���>
Za����D
p��Od���xx�7z4#�h��ehQ!�eQ7]m�U��f�A~)
�o�Y�9��8�\��2�7Uʢ+<Y��K��+"�G~��E��|�Y����cf�(Fʬfʤ��5Iz�X�|��1|� H{6D?��^y�����eD���4
d�& �.�g#�?��TK�Pk=��Q�w( ��*3s<�k/Ͱ2�!"ռL�iY����ئs��~ �(/�Wm�.ル�����d��,�\@Y���| E�!�p����6@}��kI����Y�7N�Ji�u���.�?�}�Y�+�È��U��R;�|#��?&��!�K=�AR$��=�����LxJ�����v0��D`"M�NkW��� "�L�J�Q Գ6jZ#ٽWMF�ע>[/�S�Bn���tP�A���#�����ab��`=w��E?��J?꣹�P�h�A�7_F���[Ռ��I�!��$�γ�A�詈.ss*=�@~8��Ic�=�F?���s�%Bo��Yw�aӊ����Q�
�#�an���7�RR����,�Α���q�4�v� 
�Ǖ8����4|�W�H9�����*�Kޏ�� ��R��_����c����4�I���q�!�ح��<�j��,�\3:覟�7y�o�w��a8[j��d=�b �f�A�$%��QY��g;f�@`3]�Ŧc�=_跲��%dg����xڿ��hE�8������Hѕ0��2x�g����jHX�p/�$|���6��Ys�~PLsOk���n�e�i5��DD��� ����ح|V�a)i�ܔ�a8��<��b�ފ�Y����M���h6u9�(�7'`�h�PR�;.���7�C�(3����߃%z.OQxj�?ݘj��԰&�K�LЛ%�X��Q�ٷ�L!��'�����h|�9�':�z�$�IYY�yu��Q�52�.6I۽Ny2�סA��ׅ�A��/,��7�,�B(G�5�>��*�٨�i4�d}\�G�G���D���a	T���f��X�ԻE� G�x���2#�m�yy%,�ꧢ�E��'�V���V껧6h���
^��>N��
w�*��PS�i��#3�<��}�пG�RG��n�#��(�2^׻�C(|/5L-�֘���IsX�↉��z�50�d]���qy_6򀒒�߇_���U-ݩ]�����(n����؝@ҟ�!��=c���{G
��d��k[�V8�$���y��~�d����/��P��=���(������}54R�s��F1���W������-�!)`��F�Z��j-�6�.	�K��s){3ş7��z+��PJ�U���Θ����j�Lo��hSUT$�ؕ�G�à�I\V}�
� ���#��XQE0�j��K�hr�t�(}����f����pHw���fb�.�/��>=)����~}�K_��ߏu����Z6ƿ\O�����6����З��'mB5{�D+A����kx���/�&��3���@�M��j:���i���j#���@�aS�\I �X.NP��a%;�~<s��KB"��m|G{���8FV�՛M&k?8 ,*ȠX�w��0W������ ��O�A�Ҍݛ�#q�W���i�-*�Pn�sC`���Eƈ���et�� ���\����E[;`)��1',���!�v~��aH�\����XJ2��eƬ�ɇ�������:xںEU3��{�s;���փEtq����}�bЍ�3�"�}��1�0��Ԥv��`uJ|\o��D{E�Ut�wg��5� ~6#�|}�3:�����׌��]���	J���q��aɯ�6�R�J=J�$w;�|Lլ[y�/�ώ�Q]"TO�W?�$ݕ0�m:G�C�ӕ+��@�������8
�;ZP�	��'�_��XR��Vw=���)Bѝ`FVzS� �+A>f�dَ����!�{�=F�b�˒̼4Wx=���{C����o�&� ɏ�3X/����2Ʀ�l��}t`A��~���%M����I�!�ݟO����hń��A;��c�L㸢�W�|ZP�m�e��h�>��>V���Iw�2�@��jc	}`�%�����O�![�k:�{�`5�S���<7��s���>r\�0~U�o��ly�7�C^�*��.�2ȴ&�ы��%�H~ڀ�7į�H�ۜ���\,=&�����{wW,h��2��Z��"�5 ��|%$�B��*�>�����~/ �h��U�:�F��&�c*u:��Lo��Y�s�� ��$���G�+	[���G�	P��e����D-o:&�XD87C1b��7��x�)7r��=�R*ex�a�hx�0�� |d��l!"�0� ��͉�xg�ķ8��JH����%~�p��b[~�FN�1�D�=�INo�Lީy��4���}+�����1�; [��' `BH�pe�	&�E%��F�Hc���.�-)�3��M`Xj���p	4�-"X�`a���ޓ,C�\��HmF�tW$�0^���3�e�v�i�	�"�,�6#����:ާ�A��&��tkFBbcn���6�V�i�r�;��^�oQz�e?Z��  �+���t��!plD�"G�8��
&����L7�V�����P$�7B�k5<O�m���������ZJ4��V �t�qG�Z��Wo�w�]@w�:�Y�tة�W��lxP���wc��p,�R'�X�4��ek�X��W<�)�sk�v^��yn\ԅ��[9;"_(.c!	i��9���yIʚOX��J�.���	���d�/9sEr�o%�˻�zFk��p!I�O�"�+_p�G�F��T��L��q����;@�1�h�S���tg��'u=�e�zɷ��}�^�-�������uT`Оף�8�6�[��\|�Y||��Ϳ��PS���w:�VԩF���s�Ϻ�}����q���C�^�Ft��&�U-�n��h���~�^AD���c���U�P�����;I���#c���n�Z�B�?��ciQ��]~�ٞv�u�Ց��#WO�m[J�2�R�D�	]&���t\�l�Y����'�� to_Uf�/FcldLa��#�͇a3a��~>���J�IW|��j��/{�:]d�?I���^�
��T[�
p����(�A_ e����w>'�����Rs'E8?�F	d��TK�E=��]o�M�م��QZr$��c�?1+2�6��e|��x4�xn�G��9�G�3U������Z�d�t��Sv�:$�>�!��㘖��&;/R��r���ɚ�E��{��p�:����n9#KF4Σ$�(�N��3VU
����5Z6�V�L��[6s��u����v��Z��p6j����ҏ}�%ܤ(DU3	B�c~���]z#��"�SD�ῩAe�B�������/�YXԺڇLPa�q_�Vۅ��,���s �S,��
Ղ�-�E�]��������e�rjM#K�)�^��PzW�c��𴹷�W��@�i��wmw-�C$��$%�R2�����2b��3\us.�\9��W�W��.t����+gB��̧�5�7w�V�����h�~ȓ�WЖ���،�^O���3�Ax���x���9����%f!����3lᤚ_��%����B�75)tؽ�ץlKCЙ� �{Y��h�m��bB3�o�X�(E,�/�*�7[W�@���Nd�'6�~�;D����μO7�l���`eR�T7�:�Vs;���{�3w=v��T�x��?r�)F	r�}�
؝Ϙ���n�l��M59͔�"�jAS,o_`	n%��4}*���Gjy�\��5�>Q�N��:��T�]�D�ʻ���#3}OP҆�H�b����xO�.������8��3�C'|���&�9��J5�!�D�2 �����~��T��2�����TϦˊ{哜�|�B�!��Q'.E��#M���n�d ��#;<8�����-�_8�ݡ���?6�7�5���<u��I��Ьgc�5x��O
�����q/�4yۇ`��^�^;�v�;���槨�˟H�ROB4�_3l��E���kT2�K53V��6���c���c�+S�z��y��̓�3|�8VjR΍�h}&��H���2��}���L��o��/<���".x$�`8c���䐤I�#�wP ���#�-F�)�UKN���͒�\��dxl�d���j^��E�jFQ���R�pT��3�9�p}�8
���,�m��d���(�Mn���{t�>a*�ӌ��"Ϣe�uU�P\vj=�}�^Cȇ0��u��lf-�,�A�A�6~Ԩ]Š����v���6���;�F���~)'�BO�����VyG#�z������4u�k��D��w9�Xbro�q<.���Ug��`�I�pam�!�v�*��6�uӷ)���e�c��ض�%$�*��plp�cO���������b�Ub5�'%�c�d�&�[�rO��M��4
B����A@)�*!^=����o��2L8�]�D�Q���W��������v�x����F5���4��� V�f既�q[�z�f�������	�K�QO�[0	�o�������XP~G5`��=Y�_	�ul���$��;u��X1_����Pg IXk&��p�� ��/d��:���[���A�\���K� �6#ðH�L�N��������c��!H���� ��O�\U��t"��W��!lH���ܣH�l��>��F�,�h���NL&���%��iX��j��Bs�攇������GI�u����`��n���2Q���
�����QoO
pMk:n����&=�D��!�y�0��k�x�3h�COAE��ɺ6�u���a�h��4z5�(;7�`���"�~}e$ܸ�V�����gS�U?Ո�[�����!v�t|D�ĶTìSy,X�`_֡\�������O���ȩ���^��i����,��#	QB���oʳ8��kj�>��ca����h4T�b���dn��{-M�p��w7�b��˖\�X�^B����xu�����KV.s�.�LS�A�������4�CKt��@iHw�p�8,R3�������?��R��je�k��J���N᧣��
=���d�9�������l�M5�ݣm�rÂ�aи\P�^��K���`��U<�TE�#��TJ'���#`6�q�
�d�9�]{�6�Q���S<�FwLAY�L�D�����b��������a)�87g��2�tq�L��_��X< y\�m�Piާ���#U�]���,⿇Ͷ��H��xT����T%Q�{p�;qT�$�z��tУ�t�u[ͽ�����_M���p�-Z�hS�[n�	*�q(xEp�j�#�>fW��9�0hzO��i��=�� ۷t�4�j�+U��\S����,��ׂO?]���0�Ӄjv	.ҹ�AA�����|�\�;{�,,�Rս�,�YVm�;�g�A^"|L�������7g��إ1M��?G�z�p�j�rmns�YЊf�~��Z���lL�r'�ԩ�Tzw�|��;���mЏ�-n��� ��o�W��7>PI|��l/ �2�R7l�
Oy@����yE��BPd�>5?��ʣ?���1�l�w���D��+�psT�ǈ�]�Y���X~@��᧒��V���<wI^*L��_N��וl@�臎��@R�H�p��`�:����C��������.�N�FbL�b��0҂���`8�c�l��8�;]i�-'�,��!'�"�����q	�K��{����>��0������[�/�'�PD�^�Q�s���~�vdhg����)1#S�O+�k!�،�f�dᏯ�@�Nz�Ƶ-�<pl�F���-� ��	��-��i
2.D���xC���\�SJ�ꑕp����k}Q�O��d���Zͳ�祖���q��)&�T��<j-��Dl��3� �hp���E�|e|oo��޶��}��:|"�︝�M�C4"�f��	j���J�Р�yu���6��S�B��$�ͽ�̝&�7�x�8"��%Fh։��[�Z�.�Q�pb��5FR(Mϓ���0�Ύ"r�f٨�]ȕ�s)���x���=gM�]1X��R�A�.�_״9Z�۳�"�2�B��c��}���$�U��WfK�&?�R��^k�j��@�Ѻ�d�}�`�c��,��f������g��x���,N�Х�*��/��i�P�C4Vy3z��铈�֦�n��FlZC9����7	��X�8�/��>q���"Τ��Pv�=OT��	�')�(��<1�%�e3�%@ԃ�o����Yp�f/���oV2���`+�����ͦ�R��kme!����L�j�Zz+�)��ڗ���a��3��0~0�Hw�"zʻ�²�i<o'^�+y�|gq��]�j7���_���l�vM�z���&)����<��!�J�k��R�@��a��?�&��(ƃ��φp&43 �!:s�{6���F�@�:#�dJ���7r�WgiT�
���P���]-&���H/U�Ǖԍ�$��Dg��C�G:�$ �,f���`�����ՉC]� �6u	z����5��K;��ۂ���nc�^����K���4�A(���U��5��4��^y�m�f�$�57��1.OS�H��f�F��FCE�5 !τɶ�췫��K���<�t#�Ζs���W��kľJ�L�/xn�7�*�����A��(�m�ċ�
��C
�?O+�.��j������d���s�=�"A�]8�7lHQ�X݄�b��}�_jBA�,h�6A��Q���pޝ�*P��2bl���e���<�e�Z��H������x��T��|�s��F(G��:����S��2�E^5<�s \*~
�=
`._������L�B=>7��4����V��x�(a�LU�>!2�xI4N�,8��
�����%l��Hx�OY���N���'�%_�
�s6s5�qcZ��Z�u2�h�%d ��)y���	36V��i���}әn8���B�����9�[~�Uq9q�vC����d�����o�H�̓z���G �,}h��x� �,�C,�&# �(M�F�|���X������I/�� ���E棈",�@5A�7��*��}_��}�:\U}��p���;�2��h�O-Í�PBЪ��E��TR���Ĩ�!A�
�������k�g����ى��,A�I�-/b�mz}+_sD�`n�<����bqB繟�����{&oI����kA�^K3������`�(*��+B��o���n��c�ǐ��Nj�b�������,���^�e��E�P��״��'I	^;:V�+L<�b�徵��l�G�Kb������q/N���R����OU� ���Ժ��MXQͦK�h^���Ě��y�Z�w����9c���풿����!%1�셻�Y���}��/�pb��{�0v�i.8~��d��� $ u�n,P^8�rv)��05�z��|3�D�+���t"�4���� p�ȑt��W��0��0���<�M��l)�� �x��pY��MJc�v�Z��?�u�1>"�Cޠ1���e<dF^�|BQs���4�����-K��Ϙa,-�0�jCoV�p�.�O��'Ҭ��x)k��'�X��2û�'�[�Ѕ5V3\oōiф��b���� [t�[,V|�) �3][�)B�!�S�#��G+�zv7�>95!����[?��1/��(A�r��u&��c�����/t�q�����O��j����4E��R�S+�ɘ8�`��G�_�*9�<������u�M/��كq��ҙ������/�\�"���O��8�J���ۺ��X;�u7�|�b�6���b�§NI���ə��2�*�i(������J�@ݘIƱdb�]�DM��,-�|F"�Y��,y$��B�ꞗg���#,7ܡ/��"�b�?`D���7^�$Ҳ2.���E�*��f�T5ld�y}���3�Dߒ�B��tm���W�3�`>�i
Df$���B
T��La��}u�"@�xCg@YL�����j0��Ɂ���~α��B��	���;Q�C[˓�*�Y#����YAj_IwKԗ˛Ȟ���^3Ào���~Hg�O�\�eY8ϻ�V��r]�.#�H�j;�g���Wꚲ�/�7H��L0k:#�:9N6�oPa��P�a�|砷��ScL�a�Y�}v�o�a�l��i��U۠˭�3��?"�\hFv5z�Dp����N[�w��SH��̀�8$K���������j��-=�g�lƋ���9��z����U�����D�zv?�bv����=eر�}��A�����Q��m�
GDwRͻ}Nm����{pK�����!)?1�9?RS����3A�%�g�������r����DA(b���\��㿏rڟմ&���~��Y܆�����'pC�P���D�E
??�υ��(бȃυ�5X)��/�{=��Ҥ�/3	�l�(�'w"� �'*�|�Y��^��<3����X�P)�+R8T���&3��d�u�P�FDV�e. ��?w�{X�v����%[-�C��7�=q��_	�m�|Dr��-�I=@-��'�z��\!K��ؘ����/P��.hM>�G��N"�n4XM���u?*9���S�^ފ���̈�mł7
��]_"���G���e�>{�o�oבLjrw�F���dP)��.��Hay�x��b[�Jz�W"ov�b*[Y�XqC}��(� ���(�ބ��e8�[�}~��(:g���NR������*����1�*��e8�~�QW���9/�����N��Ok�߬��*�%�Q*������=�Ɠ+���-z ���Dŧ����qz���Fё'��9>Ak���T�?��(�K�ܯ�6;I#�b ,�n�c��sp���7*�H��'�%NXN��lyn�_(y:/A1(��E���`����
1 3�~Fp\�HѾ-�ިNv)�k��m���������h��t���3}�:r`3�J��82m�R�A���lت��c'@��w޶8�g�)
����h/?9�E)4`�w7���r�`�M�.�w�8+"yh�"���&^��O��.1c:4��T�u�!�F���� x�������'��Y޳��y*�
 Oձ�;P"0\D��!	�/֑-���P](�uk�&��Ε�����7rP�,Up4��
�K#y(�(���;>���Z֥4� r��4��9��8��=$G^��	l������ؕ(CeD���Lu���@£s/zTEj���MI*$��pp�t���y��� .h�R��OK�'�_���F[X�fh.ʩs�9@�%¾��8����ڟ4��w���0}U^����m�hzj�,�c*�]L3�i�Xl@��#�]"���`,�[/p�p��OpCˍH7�C����;�^�/�d�%�atB�k��&� ���5��B���kj��ޮ�dv�gJA�}O��
]N��cPv���y���"-��.R��{՛�.���اn�����bet��Y>M��~��{����E�vs��v(;�t���[)4aZ��j�"��1��cUp�TG��{���r�\���������������Ҝ�2D&5���_�'EQ<�-mu�΄��ZuFj0<\�Ҷ����nkq�A
�	�(U�3L��Ȗ�1�?;�g
��@Т��2�~.Ƕҙ�����d+c2����J�'b����o�@9������|�TL����y_����l�!+�B�Mu!g�=�Q�0O��Q���C�GFBΤ�t���dǂ�����٤�֘bZ-���os�B��L�` L�X��b&*Ռ��[(7� Z�<�0�Q9��@ƅd)t:r�^�����|�&G���t�eI���g����?�#uO�H���u>`��Ls�K8��!$�q�(c6��W��z]s%w�y�Υj��;tR�h��ee�oVA�M�gR<DҦ���^>G'bC�����8�X"��S�F�NqB!0UngF���-�%fγ�+���iRtsϵ�90�!�^�^4�o��]����4,S�xX�����[E��r��B�A]	p�f�|g�Eu�#.��e���=~Ab)���Q��. ����WXܽ&���U�t�Es�+'o�f��*qcb����C���3�8P�oka�P�g��U��&]��1���`�����MۍJ�I��ߝ�'��2�6�`��'F��lRP�^�1l[6Fvr���'�E�b�)? �a�\xgK��ɰ���pE��� $�£I�{��У�.WM�i���~����7��h��J�/���Tp��<���I{G 9|76�)c��Lo�i(lH}% ]��j;�a|<˃jQ;<�@1פ�t�+�T�O|Z.��+>�ًu�;2�ȨL�_������]j^����ۅϤ���c�KƏ��Q�@şzӄ�|�܋�W?h�� ��ESE9z#T1=dժ��+9��D�[/ݥ��z�{�6��FGX�Y9gEQ҉�'G�ӳf�s~���?7��^L6�z*(�w&�*кu�fmR�_��	�[J����G�`%/N5j���ӄ	�e�O�ٽ�bf�GbQ���2�'��u��s�Bg�p)�=��B�������)ֽ؋��hrʐd��L�,u�O8�2��rKǪ����ַ���9�_i�;P�u���P�d����S�|�~ Ig��Y�x�i��>l��M#� ��4ƥ~s5���g�5��=z.�.Ѳ��p��٥H3$L����5fqr��X���B.�	A���9�@�=U���Xa�L��A~���%��-���侍���:)��e|?>m6�CŜ57��A���y1���V
�D��̖�U^Ѻ?;�g�fN�g��/�,R\x�j�r�����A�K�k^K�5�r�Z���� �4>'����n��^����+�{Yu�5ۊ�`�:�1R�As��{\���!�df�<;�C���=l�hT	�����h�T_��7��$ �	���>�k�g��0 %�	�B+W��" ٍ���mV�z�����=�\D�g��s�Wӣ�O�ZC�Ҙ��ckJR0P/�*��pҙAo��ʃ弙^�Z���e����,���j�_�]��EZ�`�_aI������Z&qi�4��$�t=ٚ '��8~�M¦��.��e*�P�*�<��B�E��p�ۨ ����ʀ�h��_W��s����?������c��~{I�j(�vG��� �����6�R�7�/ƛ��HC>��11ހ��ς̏���MXmΖm�i������$�}<cq�/r��E_�}���"7(���*%�"�k�%���X�K�R��d/?Z��3���A`4+�`]��N1����T*J��y���[�Z��@���!Y?ε����ڄ�S���'�$�`X��ŭ�xCpC����)J#.<�f�t8�K��|N{%\�����{9��+�k���x�_8�r�����B Iɳ����EG;�hb����	�����^|��8R��*5�� �1vA�����Mb��br-"����8וN:��V������TdLC���
|2���N̼f�H5B�\��dTq�����(�L?��|H��(�x�"�x����$�����ͺ��,ݡ|�-^éF�aM��Y�����cH+��
��L���,�A���_����ع�:���P����[>�u���S��[��A�B]g���إ��RFD����,$�����3dQ�S��R
0��� HL)H��Q�r�63n��t}�Z�RآO���<�٥0��nd<q��w"�[��y�!mX���]�1=	{|���o��(��20�lm�yY�s�ׇ�C�\��ў>0�[�uo�N̗Hݡ��2"�3�ح;pq��;g��i�3��;��I��^[Ȟ����יBp\A �5��u2��{la��Ob���'�dס*x�Ħ��N\��g�P�f)�E����d[a� �3C�G#+{�W�ꑂ)?�	�g��������j�9����y	�+�����[��I��5���B�ӫ$R�����&>����T̂�X�I8 ��oR�]~V��[{Q{�7WbSY_oim���3��AqjW���MXd���&o��K�����1����21>S���Hl�.�B���%p�c?ir�U�k�����"���?�rn�����;���������\4���<ԑ��G`���A�=dJ�v�xY+"�}�O*�z�������ٙd ��ˆ���}�@���g���eB7�!�e�:��j���rwAY�:�XO-��Zb��oo2�Lα�} �G9ǚ��j��l��w%�*'�7�Y�z�xS��줶���v
�A9 �q\O��y,�A�j�H�$_��h��tl sAГ7�:��&W�<�W5I��~/a/�rųܤ���&g���J�	0���ͬ�cO�l	����S>�J��֫�����U�>������`ҹ[wڢ�^S�V�ܝj��} O����A�Ήc�*����fPu5ͭ�"�!bB�Z(�vUѣų�.dsמ���g���i��yY�P=�W?�nVNp��w`�P@����Jvڳ�Q�9�HI���*�c���q�}�W'-OC�R��<v��N�45WW���>[(��pxUb�t! r@`r�Ɏ���ъ����=0�'5��`�v|�lgs�_��x(,��|������M�{�P���|�(BL��[�	r��#�/�\��rO�T���`V�/�����䃴�c>n�I[fӤ������y&-��7~�i���`IL�ꚝC�ϓ��}��s?���$s����F)�kh�+��$�Xq���DS�$b�H��i� �o����#^$F��uF����d������7o�/�ሲ@.���~9����F�����hx��Dx����s��c��k-4Mń�W)�*���b��s��@5���F��h�(��$��:����۞lM�]�c������UG��"��oSA�c�^4���>"uΧE5d���A#�f���݅7�m�9n�%=�ͦw�%�H<�j�V��cB��Z������hS�� �d��;9fy"ZMܘl8�%!|eX��Η������ �A#nр�:2�ʋ���ui��
�ƉU��2S�:����V��9�j3=��'��Tq�I=Ήا�d�� �f�T�Et{}�a DWT� ��cǔr�[�f�QQ����<�E���V:u����Zi���`���^z� �|��4���W^��);z�Z��(f:��P�,�Q��>tCƁ��p�Q���Q-ó�!!�<�{=�Ĝi5f��y*0�ų�C��V��l�so�6LK/�ƅ|�Y�v�+��?�#�U̡�䋵���2�C�͊�C�	���݃@j����F�!�^��r(50T�%�
��ta�P��}k~Fs��x�]����a��(�zd!�9l>.[>buM�=�=�{N%f�o��~�y�_h(�gMq��8�8P�Biv��Ok`'g 5��4�v�������;~'��B�=d<ϴ8d�|����tV6.����@��V|Ɵ��S��e�q��QF���b�~��,�8
�+��Oz|K\LDz���.l��!��.���IT��]���+�_�jiC�����A��~[�c^Xv��� �Z���\T;6uK�Wۈ���@≓ll��Ͼ�rB�����)<�5�����Md���t��SY��[�Vߨ�Bn���wm0�]U� P�����X��4)�\=���8�#��<�ģ�E��,����B�=�;���/�ٍU;)�Ѭ�日�
P�a3����@f��N��dT�q�S�w�	.�	N7����]W
�'��hY#f?�;��Гj)Q�1o�S��%����*��;��iچb3:y�tM@�>�,�d[<%wt��; ��t�m0i�H��O�~����m�m�A^��.b��Y�p �gl*��NU�D/��H�e��"��I�f��4�=�Ϙ-��n�z@���N��:��X��ѓ��p��/��芴�Y����❓ _zBe"�4��Z���
\��8�i᮪�=��b�@�I�P
�����ȃ}M��v�&�1��z ���<ئ +N��K�<�̐Y�1��8o2K�	6���b�����g������B1�1W�7�X��]&sG'-J9��m
�ɢG~��j�eJc�Vp�'��KR}���V��6著(�А�iP-�m�fz�:,���_ona4qC@�4�{Խ�ͩ�<�QܛA��c�eWR��TFb4^��K�Y
kdF�ڳ�U�)��[�Q:F�{�ջ�1�@p��	�s�;�H��ne<U����D���Ȩ�V_�X���tD~u�v��vV?������-r9+�x��;�	m%��}���h#~l(����#\�jC��s�3�
{��Wi�E�a!���Tg}��T�*#�{dRG��7a��+s��ީC�Nn�C���"���"�ƛu�=ٌr�0�.9�Ì�"����*��_�tN�8���:-v(��|����Ѷ,�d%�ѴU�
=�y^iwOԝ�7��EE�6R?Uz�Ӟ6�v��O�M����qa�$גw>�/)��E���8E�}���U�tЩ��OsmfQ��E�"���Z��ӑ�
�Œ�j�@}��l^{ۗz}.4�3�%���7�q��"�f5��s�w�l#��,����n��e.�D��l�3쨃#Nⲣn19�zW��3�ǘ>�8�
۰���<�W"^+��.�b���֚@l*Hǔ�ASl��05	��˅���eQ�2�.� ���J��<7����bg^C/
>����A9OS��A�͞s>Zb����[f�6B$�>{{'�[�B��ZL_zV_h�Ǿ>��ب�I�⯎3f��p!"8�N��_L�d�ͯ�؄`I�5-�dX*���{��N;��[W�>QT��`������~T���L���Z�z=.���S
eL�d���z�%�����}eMnF�볲G�d�]���&؜}��������Y����ʭ!Y�1b]��^���#��V�����7_>�m�ΊA%����i��-�bB����<��7��E��q�3�4dd�{�z��"�j��^G�^D~��kQ�d��!�zD���bƣ��;�c�������؉S�s@f��lbB�:6]M�&��Z��f��M�m캙S���1i�_�����1��V�5�HQE���O�� ��pS�*���st�Ț�Om�TL�</Z�1���U��r����U[~�:I�	o�%��V��Y��=u���z�氘\y��b�t�-r�p����۴
L`�	� ˹aRL�;\�F��;i�s�ZP�Q���ܭQ����t�^��V����G��<�.�S��)M^ܱZKޘ��D�g1-�������m?��=ң�G���8�FM3��-���V�4o��ڌ��T���U���:��E\7���#�Bg�7X��,���Tl5�ϴ�T>�	8���D�3�r<oź$�@9��������0�>4��,�P�:��9���8��X���Q"h����ջ�ߊ�j'��|��e���*��c@ E�<(Qunw"? ����|�:G�G��Xܶ=�=׸/��F�g��%��?�F�-��d�w�q��9�`j�� �sk��L(�3��/�-�o�i�iZ��(Q�ۖNt�� 
�6S�oN���l�&72yzT�b��{�\��v �ǆ�2`ҞˏX^ݓMl���N�o�l���P�@�]�O�Py��t;�Z�#Z?�{;��bHE��ω��u��ۡ.0e"��q� l��	�`�T�r��t��^�$@/��8SDGе0�`�e-y ��\�5���n����0�N���כi ����I������d���Ȏ�F�B��v�J@&�߂��ܟ���(��z���F!1rw<]d�X�c�c�|O�}��X���;
N��9�B~�F4��<�pHC� nҲ�xI���وe���	�bN�]u7}A��1����/��n��(⿸|8�#br��$����a����ޗB����+��J҉y�	>��2?�n/�bVI93t߽)�P�G��0�QO�%'+�:9e��Ne ���@�m9RW�Vc���%�P���p�&�M�u�;%���s�����ìq���z���������)5����3�x� ������`�ܮ�L�t
>��&��r6&˗_B`��a�s�.�]F�l�v X��(n���j|#����@�۽��L� �a�[��v�B�L��p�zN�	��<�&��n����?-�E�jD�4oF��_ �� �LÊ����f�*T@�����o>L��aMĕ�����w.�&�S�9�����Ҽ�v8[�y]��J��i�&*54)��4(�q���r&��uKOzZ�[a�(�F�� �'S����Zܻ�tG�+�H@u%�K�����N����w�\�SE�J�<Df8���{�����U��VA'���R��Wo'�,)J�,:��.�K0�˼�'
}*�p�$�E�	F�Zb�qŻ�)��Af�?7��@C=�[o����a�Us��rMp�wf.
8&��_8�NGEp��N�d_T��-�"S�R�["�?�%P �c��x �}���� /���	����Y	>Ji=�LqUF�of0��F���p���y�P�ѕsg��/l����H/���>��I:?EC���V`Ц�9�<�+z]p�-v�"�!�}�|�L&�U�'�-�)L��S�4O��~��Aq0Vd�o�u��Op�oyP��$c����ڊ��?��&js�g��|�q��̅by��(��Tk��w��NT(�q׼H8��I�"7��ZYi��Ԗҡ/�_��L�)�&�>#s�8�L����R�R��?���_Q���Lq�!�e����c��� e��2r�S�s^:/���N*2(�R`'6�:�ų�>�|�G۳�s	�W�LGX���ɀ��H���J��R2�k��'��˞ �}��?���n�g7�U��f1��N6@ᕔ��(+j:��l"4����<�-�U��G�uAXt�;�G��Z6�A�]�06�����~�)�w��	ҷ8V�����z
�}F):Q��4�6�V�C�S5�z�ʮ�)d!w� ��`�'z��>=�����`r�8Mۡ��G!�9�3��M�t�/1}J�ץ�L��z��7W�[��{�?[�y;��T6��}�-��p{f�m|�KZe� �<c��c�[̘h���MAƵ�`p�a��n37%1Ś���������������6���nM�_X݋C����V��wFa�bo����)ٽ"3+�b�i���U�[
�g�a���42�J*�@��ۍ(�Ӟ���>u(���r�ä���u���-NяX���fO+V�sEv2���I�WS�ݭ3������H�1�Uk����݇�(�8k e#��7ȃMAG��L�S�X�$�1��nJ��fBW�$I�rR��y3(a�أ���,$r�ʪ��-��qK"%���T_1h==����lǻȠ��N�����ѫl�ݸ`x� ��,�B֥́�$p�RT��_ܠi�"|��/bݷ	��~S��V�s�9�=[8(��j��n)E���	�s=
��T����X��j�C�X��M���
XSs�'y-�3�iX�P���ĵ]��)����	���3��g�{�@�#�[��#�z^�nmF�4-�V�bD\)��f�vѰ���#'��.��� Y����lB�2�>|a�U<Ic��DO�Y.J��|ީ2�����̓p���o���O��ؘް���bf���؇�j�E�r��D��R@��a��t*~;e�����S���:�5�8�=�DK���U'�;�/� ���8�_	)�ń�2M���N�o���4�����8�*>5�����\[}��r��=(��*�S/B��/����%�܍�$ȓ*p<
�K-�$ql��H09��ߘ�\��!ji��WQ��f��܋�_��JΖ����i�G�&B\������1���e�tj�o����iz�l(�e�w�����w����H��>O�qa��a�,]u�{�Ҫek�a1��}�m�7��!a _��c�u	��m}�:RS*Ç����TF�<\#�������b�� �a��쾧�VM�6�>^���t{,c"�=��� ����A�IY�z/���?�E@��Du��8r�`�rE*),��E�~��6_&��a�h�Oh�AM�,V�0����=�Z�g�U�\���a�~aj�kr0^�c�\�O�Bm�;f�"l�0w�^���U��zP�b�@\���l�V�<���
g����E����%��3��G�5D�wg[  L���?�����^��}�zA�sv,�F8�F�5s�x�LD�+8��|;&7,������;���#�ء+�.�w�N�N(.b�w|���XB�Ǻ����ؔ@=��ou�'�3�{'�4s�7d�PB_�M� �XJ�i4}��'/�T���t�1nw�,3�b�:m��ْ?�Q_q��/�B���_�MWN>-I��1�@�J�+��h�:�J���9�c�U0�qY��%%�Ϋ��р�1
��8�<|(�W��W��*�B���p,���:��w��U�ILP�/�ʎ?	�.���c�n��Ɣʃ4?�}��B������T,c�M�[�29�e�f�"��p�j��5���t��#����^��b�Jy�7CrPٿ'��8ueҙ��u��!�^���}Fͼ�� B+�j��GyJŮ�@���".�0�W�@�BH��ܩ�]{����\*�W\���Lo��^��q����L̓Qۀ�UQ�y�����r��2���dǾl���&�Q1����,�G]G��v�9�$������(Q� KWU^ޟF5ˁ��v�~~����'�Y��5�U�����;�ۍ5Q���q�b������[��T���b�wB���1td͛��D
pĦ�)��֪Fd�fLrWAHj���:�[���Bi�<��+���N��Kz$C��;E�.�x{����i&�X��˨��l4[�H�
�H��;:�:�m~�?�Ļl0����{�_�|(D��@����BH��qa�1ˠ���Q�[�{��d�N��N"����/HI��쳾��sg�M	��mIY'0y��0�<�}�{��]��;�6��1�yя���D�_zߘ-m�Ӆ�)mV]��f����=�~��1����9^'��=��ae�&>[:�'�I��<&�+_Ktf%�r��Nkꑼ:<J+ǥ����F;�Y����BxlG�yE�7
.�V
�Í;B	���o))#�u"�,4���M�5�NJ5~tk���'��ij��8=��huM������x�]�]A��6�����yo.`���_�X��|Met;��<S&:v��-�l~az��I������_��+��t��k�O�ELR,0/��: ��_�Q�V�;v�w;1�z\Z\�e�ƴc}��-�	e_�+�x�Rъ���1�z��ו���߆Ԉ��?s�Q>x�h����A�w����/�h�
;��� �J?;�.�c�%>�)����I���H���P@2�Q��_��·�V06%����K��o2.:2[�/7�*,g^I�,]�pO��S���x��Z����j��1J��D�c}C�.�����6��y����]��f^8/ o��� ܛ��o�fK��.U��$K�4�X2P��=�]A��\�S����g¸O'�fV#u�g���#�+��A����A����� =s?��I:�a�Aر�B��у���=���� n�l��ւ�Ҫ�HE��S���� ��˴8D1�}T-�C�6��DI{'��k��4�S�|��p�KËG�*���Jѷ��'�.	Ƕ���Y;N��3�@�
��T��c�^�9�	�1p��i@'|ӵ�}C�0�˘�3�<��K	�TK�i���&��{� ��&�b��o�Zxx���Bl�A/5�s+�BpB�2�l�?6t	2��3o��S���I:�p�L��&��i1�'��bY��s�?�kq8D�Q��v��S/̤X9>ڬ ��g�)�N�l�0���	��(b�8�`V�S�cLWe{p���
Sg�@�� 9�����m����T��$�� KQϷ�$u�g��9$dX�gP���wU먂~��tT�G�����%��0]d�H�:3j^������\HsX6��L�j()��v'�/��C�a`�e4��ߠ�Xk�t#$
�Ɏ�!|I���'�;�>��;>�����0֋g���~�BY�ƀ�ו�ծ)�ڱ������C�I�e��Z31�o��=w�80�g�lIv�_{m��JSkoՄ_����]��W�%�'a��1�;�{��!N���F���L���?�zn9		�&����7�0ň��V�����7��٢�YTG�Bf/�&-j><	�-y6�6,b�T�Y8�w8����4D�=}����I<����s��^����ړ|:rץ !��9E��L
�s�����&�R�?A��֭�rko�E��&�ܼ� � u��y�@[n�^�(GUs�n4^��e ^��f��I�l���s���F�Éܩ`�Y�R�jg�&�Ҵɐ�@G4�TS�5��VB:`�}مIЂ� ~z��]�eF�Ѻ�|������>���,`��5>����ѡ���?�,Y�m�8��i`_X-�A9<��
�"�jyQƆ��y�;�C�����VJ�����Z�a�[#�0fܣ�5w5 ޞ��>��'`V�ȘS�/�,Q|��CY�q �@�8x���@���~�65|��V�Y�"��fu2+���� �:$���Zp����*��%Mq��UK�GIHW�5t[��ݤ���#��2ß�}�R�Hq�ձ�C7ʓ�D��0��\��QW�@+���(�,���m��_��
�k�IMg��M��	��@����#X�k���2��L���ac�pHv�Le��]OIs�iu��	8E5�O�vzD�L���`�u���$�i(dSܐ���*f��ɛ�u�l3m�U~��2E��2R�~7�qi�hd�{?���ܺQ����ܠ����FP)��f�5�5��Q	���>[���nps$�Iq�2�Q���( 1]��� ����튣���xu�WɎĐbF�
OM8�PZ�� m!�4�x*�%�0�錍t��U�����p�	�@Y�Gv�ɰh}<�ԃ^���h��q��`��>���a�o#�����P�Bq[|��%�a;^@����+J�Rw�J�ffj{��^�X֕NQћ��}�$g1�К��h��@S��q��H!�"�b�PO0>�,:J�������E:��%-������)�+�*�۶��� F�
�Q{��0�ڊ�ք	&71��r�f&ߗ��
��(���v��6)�;Yg����-�_:b:\n��c���5�Fz*���������7p���i�bJ�j:��f� �g4|�l����:A��֦��_n��s�}Z�	�����[�v-;O�� ������BQ�6<��|����E����g�g���p$ra��8&��1� �A��:I�m[F�;�1�����c�����FF[\(a9CN�?���-��?X��9t`G+�*�Jcr���oJkq>���Լ�k��1dV�+��[���=
a�v�u<��*xt05eB�����O��֯�W�Ox����5?ˌ�b�xSR0�e"�ȵ��[q ����H�۝.υ�P\X��VȜ�~t�4�客�%�����W��UH�m�O]��~��/;mJi������'cȀ�1��+�`a�Xɓ���Z����E?lo��Գ��Au�!�=�.oT��>�[�����i��u�R�3t��K�!RŐ�9ךB��yH�
*:���V�޸�������̹؀�Pj����]/������X��X�~��e|EԱ�9�u�VA����t�g�T�:� ���o���Ύ���g^�L��j;�?��R�[3�ãb]А�o��J{�J@V�Vx�[�:����	<��AZDH`�e�BDVu~��f<��2\���ś%�k��k�H�I���筐�(咗=��UH�%����f�0����Z��i���Ϩ�p��a���~FC�I�	eA-�������ҟ���R0FZ:�(�Aj4���v��c������Q���MO�O��?~��<�W��{,��^;E埧p l�Ϛ�m�L��m^bfYeإ#|tm�������_w���طg�]��Qw-N��nh�W`4����Y4�!����أ��B�ҹs�譬�ƽ�q�����dYV����q;�?������f�U�N<���,�V�6��\�$< ��97H���4Q|��X�5�Qm����K����<��v|�<�k�a�B�0�#f��C�>���n��*j��F�ɚ�1S�1m���`i��*��_e����#��ww��G��8�pY����)�W��M� ��x_���R�W(� Y�����it���P����Z ��)��~!멮q�뻄=�� �)��V�k���/�#I�<��d'��Y)�o�����'4�n���/;�o C�����Իf9RF���_��c͒�S��a
0b�`#ڄ[�wSO��T���6ֵ����6��'�3yl���������y�t�$獇�c��L��hs0����L��8D�LD�Q�zzT�tR<�o*	c��0xnsruq��}>�@3��^YLt7$�]wo:�gl���Z^����25n�E��7yT!�>��+wC?*G:��։�xd����|k~�l*��-�h' P�EG�6ȩ�o6��W�3H��Հi��w����z�	�^��F��C�Y������ƌ3��zާ�����\:�����~oY���������b�I\ak��)���3�e*G���A>�:JP�9�P�3�|4�k��!f �
 d�TG�d�U��¯��M��?'m�:A�z:�s3E[��@��ll1{�#�S��J/J����v�Y&���!-�+c3�Ъ�Ҫ=�\�L���
pol�CY��7;ǂ��u�5�Bu���L����3=��J}W����L�٩9�N�\��V�Q���y6��|������D�y�^������ߵ/v��l���"�|3@�?������D�
�聬��un��:���7�Ο�u�(���z���sz�A��i��_��J�l���UȮ�tɭ4���I�:�I�R*��eq4K�����p�"��ڠ�5�OQ9�s���4�p��L���@u��USK����oә3�	sA(-�o�7Pzk`Hes���"�f6gUQ� �ݧ�ػS��pӃT���yGl,�<%�&6[4T�pՇ>p�0(7l;;?���r%u"��H���ۋ��f4����
�WoP�:eA��	n>��R�ܻ�|�U�*�`2A�pX�O|��$Jn��
�RH+��u[r�8�1BJ"\�ܾ��ƈ"^c8��6TZ���Ȯ*=����YTS»�q���R��g_��pfSs�ɞ�^{MxZ����#'���J�gs}7_{
镍�t��g��g�U��VT4��d�]S�M䭝,��#�S���*D�b�¢�Ʀ^�Ʋ�����	u�l�I?K��.γ�c��ܞ`L�����k35�Cjy�|��'`���HQ�o�JOx������7p������:h��:޳T�)�ߐ��a3���?�����t��r ?	�A/8@���ݥ�-�G��ڎ��0׬aXZ�uJ����k��Q<U;y7c<g����~L3����,k�:���tsXk�/���Ѳ;ܾsć#���������`����H$�-����������:�g�z�Y�ۗ6;�Xo�@grx�+�~�j���5YI0�e1����,�g!z��Wl�B�$��l��[Z;������:0P���k���VB��d���D@�|�WI��x%����@ƕ�tׇ��f�
�h@|�09���W��U|��x��q+h�a�a��0G�ڲ\� ��!�����Z�aU���᎛��%7���M=E���
��H"�w¥jw�mF^�F���9Y_�#�X?JZ`zl��ctECg��������V�0�F=E�0�V$�>�2�[��@L��x�,������rz��.�<�ѯa ��ׯ��KNQ?��S>Ր3�Z9w��R�?��#A�`Mz�>�����<Q~�w���1�v$;��חA�8Q��v'Ӑ�����30��"����G]˻R4��]Z�!~���s���)�%p�F��Xt_0�4�ӦOeÏVh�v9���\x����J_2-y�p̡}MlH���oH��D�.�JY�2Wڮ�z1�4�*��[e�@��i�^�zS�M8~���;*d��v�0�# ���%��2D�Ɯ���!I�j�޹ �A|,@_Z?v,�d	i�ɺ��p�쇗>8~�A >_'�ӧS,7`%���y�����mw����h����+�H�⚸��}|������m� `���jN�ҳ�	�h��Fa(O4�������s:LLz��r���K�����0]	a@S_�/�7�LN}�oB��%V����lJ�~~-&�	�a�>(�#��M�r�7}n# �-	dHb?��,Q+��1E�[�B✆�T��sxA'���cu�0h$�vˬZ7]8I�-��:bB"�y4��LP�U�����d�\Ig=����na���x-�/< I�;7�����:�K�;��1Ƭ�sМ�3��{��c�7��ͽ�:���s�tW� ���C_®�+I���U?�&�d��z�H	-����N�w�Fr慞����vL� ��ӧ�3�#�0Eu�xM�y�x��d.�*�P�+�t�kVl޼'�q���<=��kUd_?x`�a��(�5��Lބ����
�}���/�H�%�
���.^ԩ����AK��W�ټ�����)TP��D��1Bڈ3����s�#�%AA��Q�,H�_.�>#��ȧ_�r�|�c�p(� ]�Z�8e��s���f��AJ3�Z�;O ���z_"1��Φ�y!�H�a}u�=G�d���%���۲��W���߽�>s\�C��ޭN���`]�h��s�P��hP,h�s�y3��D��&�S�7N;
J��]�u��"<pp(L�Uj�S�>�O{�]Ճ�'MC��z5=��X�P�<Y��w�gO���x�����YcČң9ɰ��}�����Nܖ�pc�����jQ�i�v��<�5��n�����!����@����g�y����=;���j��Թ2�D�\����	��m�+�V��r�R9uD�<�P�LČ��s���bf��<�:��|��#��y�����zƴ��1ON΄ ӰtQ8�i�RDJc��V�hW�ݣ�2������j�}S�C�E�p\.oci1�#]����s3\�I���,���<tH���.m�n�	����&?�7�Cy+�q��/܏J�p�n�Fv��X>�Ƿ�y�@u��0��|Ǩ:�3��]����覎A�x��b�C���C�����W-�ϖ=������ϲa$l4�x���Вiҭ�K��қ��<�����/�no
��O92���.��^��yu�iQ�'YB�������4_+�ř��6��^����5x�iB�+?)�d4�*������;���D�;f�!���0�r�yc�.YmL���~�VU���J��q`��F�ҮSchB���*���J?�����ji|������J�VQ�~w�@�k*b�D�T|<�'�����ౝ�j$�t,*}V�.I\�Z�=�S���s����/@���.5=[�z/R�������0$C���X�!B�06�����x����cF\E�"�{�p��-"����?)�B�$��c�q��{�)M$� %���/��C�ű9��W�:� �vr��W(4ma��{�_���1vl�܃��A`�UR��-�[��ݎ	M.ts�R���M��B	C�����{9M�hZ��Ψ�+�����H����BJj5]��l�RN���Hf���M`�P9��M��R:���w�t��]��hU��9s��֭�Ӭ��t&*
�M/�-.6���� /��H���?��x���V����?�7*=�ƞ�:�zŨL��dH���~P�p�1�����#��2�21�%��y�]ED�p�ݬ\�I�EL0��4��|*03��~�����]�6E2i��+��M�x%�bJ
�>|��|?����c$%X�-�=�v:ǚ����j�Ң�w��F�>� ���#��(�+�ہ�����Y���5��Hf�v�0���z5?3�e����	�֞y�nL�&QXU��q�|�8���B?���}���B��#w����9�,[C�U�� O��Uq����s�[�B!ۃIX&M9���f+a0$�~H���4_�M�[�-^�O3U��WRl+4 �@rvg�H��* �o��L�#'Y�"��7�Y��'�X-pI7]��ׅ<BW�QJuw� ���� p�_� Sd�Gt�r@Pr� T�?��$kV���a@��}�� "r�;�-|53��ăs��p|��>m���"LR�N'�ǋIw24��b�\�rW,��d`��J�I��x���U�X��U���˶da�6ϔa
����.���E��l~�)L�t�d��l�ֹ��Ϳ5D۞aF,�K���܌�^c�S�f.�\v�7�'�s�:���Q��y��v�x�ʏW�_��4z�}e:u���z���b�9�N��}x�{GTzbu���dݓ9*d.e_�w=��XyRF=�O; ��,��Z��ЏJ+[(�VÕߊC'u0�IPǀ1�.|����D��׎��"=?��[@Q>x	Y���}��&h5���R0����hB�Ӯ��MLC1;������6A�yL��Z��Ӿ��.N�-8�Fz�f���"�a�t�t
t�ɏ]cU�� �����v�萴��2�Ug����N�f�;ޱy���=elҾ��є�����-�a��}���(-�غ�>Q )v�q䆆�]�#���^�1S������G��\������;�C��b A��^I6�k���A<�����͘���A���  �i��O���<{D�Ri��s/ �N��W&�f�Z�;��$��4�����d�����n{�_�<73�08�O. ���u�']`IG�8�hp�J�m�w�#�CK�N_qi�����[�"��l'~V�w\;9.�"*7Ͷ�Q�FP�RZD���tZUA�\����=`���SK �5<"�s�W��5���-ޫ� e�����|=Ai��2����*��+V �h�WZM$=%�l�v%f��4���]�Z��Q&�ݓ�#޻�[?ie�_VD��3�FI�����yXDU���1 ˸��0D����C��3)��E-���f�]Жo�`�mG����*�� @�i�*JH�נ��Z��6���Hg)mD�i�U<l+%���Φ2��]G����y�.h�tq��[Ջ|�+� ��_��]����ײ�<��ֺ󧷸��vˣ����Kj
�������1fu�<��/���/��'�7���pb�� ����P��� *�p9!9��Y5�5,}��"�{�f,�*Hj�gz�Xa�a9d*ʣ�łN�3q��R���'���n�29X�9�ں�.A%�佚N�ǅ�w��L�70�x[�X-�eȖ|��Z����R��>C,���'8�Y�5��́�MT���;�Q'C!VξAL/`�ySk�.G�M�7[�pܟ��뤈Z�({�kٜ�}�l��"+H2$He��^����.��<��)�рX増�ϟ�O��;hd-Uݺ��������\r��~OI��� �����g�ĭ�Zlb��XO�ȟ;Q�H������+�l���� j�c<+=zǪ�{mx�7�H���C]w�F��ޕ��M�J_���A��+h�Fa�;A��	
# �'MV����.���E�M��!kCl��&y�!��0�fXAQ4�BWK���F��N��O ���y�.Oj�,�A�XA5p(���\(J���Ga������ ��+[߂g;�N�L�L ��4A�ԴFU^0��Tu����}<��y���g�U����j�H�\{��@������Z.��
%3��Ӌ��"����K��s퓳�`�/$r�S���Q�;8��@����*�"[���F�Ԋ�ν�gU�07����%�0�#���X�"&��4��G5�Hd�d�gZ!��N5�������ݙ�q�2&��Z�A�Acɥ,;�����3R
�h�g�l��5Ur�$��`3$���l�S�*>��8/!?o~�?�p�:�;B���^�S�PAB鱻�������i�+B����/r�X������3*��k�fx�Tf]�l��#�{w�:RI�J|�m�I�+�*�U�sr0w���xU��K+x���y� /��y=Iŷ�n�QJ���Q2p��_�Fſ���Hx���c�e�cw��[Dŝ�2���r1$��#�AD�A��B����OIw}�/��xU�ڋ��|q$�9�Cc6fFܻ\�up�W�o�f9����7�'�{���>���V���+��Z�7&du!+֕�f���E�$H�h�K�R���Y�vzw���cߜ\_��g�0/L�|�u58��~#�����{�B���^?[�������O⿭�j7��-	�,�� k���bhd[�DITKո��#G'���#�H��02B;�=�9��yErV��)��E~R7�͍|Z�v���qW@��
XM���<>���J�_d֒޻$�˃u9<{�O%y���쐇�A��R^&�5����?�������K�4j�`-�B�U���s ߨ���.��`���Z�K��ql���oDa%z�öM�9�s,�	����"B�w���7)0*)��pBE�� �s'����PL*y�#!y����Wk����pd��b�e���f�gEP�V`�X3�M�9
�Avs��_$�`�=�}��=�� ̤�!�z�k��r�d�Q��*�4s�,|�[�z��rG1� �$��v4|2.���vYx��*�_�1!|C���.�\ߓ\��������6'݃�+�Tg8����J{p"۩��.��Ď�Ѭ���jV�ɓ�\
<�:n #Ā��J��?T���y����{9��(���@V4��G�W'ѹ#QI}r�B�ɖ�����zgY�M�Yz�[,�hK}�T�[�*F�c�����k�r4�™�Tg\�$�9�t����,��2e$�b蓓��%�j�ﶹ����ٿ "�n�k]�a��e��7�0��o�5�j݂���>�z�zH���KM�1W��p��q���ݨ�Rwȳ �i��3���65���O��mT�	����~��	�x'\�9�7Y�$S���7������1H�/�����5'(E�}�&W��n.��-�-o�h�8%��2Z��Gu�M�V�*]�}i�ɚ�ӽU@�Ws�G��R.,?��-��f$�KjEc�Ru��w+S�,\��(���˛�LP�I���-�ݩFQ�X���9l��S�+=��Sw�%B�t�����JN�]m�;?�7ICPD6m����� �B*��;����|n�M]Eb�r6�b�Q�|T3��d�#^���V�P��p� X�'��RR�\����/��� G( ����5sh��b����]���f�E�"�;~��o^�2#����''Y�c�yǉL��^'�zAILt�	��-��|BS>�!_=�8ik�l9��7�c�OP=�tjΚPbݪ�����ͼ�&���<��\����t�h�C��F�W'^an�e?�͹���ϸ�Ն�n��O調������;�̍T`�x�i\W���ˮewC���a����k[�gB'Q�0�,w0��k�;��n�Ϣ ش�g�[�t��):3�����&����ރ�Tg�z�q�K3�!3��hZ���?@�y,d�;U�K�^�ydm����<@^�PO� XE����������!�E=u<�9�Ӳ�CF�8���}=�^�O&)�������b��|K���ȃSQ��P�ݴ� ����j�A{â�v�2l���~�z��$��T!�^���<ej�������q�TzG^�{�΢A��XJ�?6�}P0<�7 ��ؿ<��w���Omf�6}E�:��$��nd��}�%���+f�Ce�q�^s��5�9��K��?{<�PUY��:5&�o03�Zq`;��M���L�#J*/�f�
��#i�	����z���D��:q0z�ʞ��Vۢy��k�����)��a��թ���Y�Ǟڸ �$�f#��yH8ͅI�Qj��=
�ӝ�ys��DZ��޳���Nv`�`@2���? �I��2�a�/��1=l�I)�F'zYZƌ75Ӫ��n	#��7I�m�Kq�I�Y%�J���V1������P���"���n�%�e��_��h҇w��ŉ���Kg�9\�:���]RuL\Q��K���;�E�0B֓:��[6`"�ԣ$>j�S���J�Fr�ɩ���#����=袼Ǿ,V�ӫ�Ȏ�m�:�9|�dRI`o�� @����N��b	(%E܌�?sdP���������#�1���8=͈^��V�6<����sopwҎǤ�e�q��FE���)'x�ɊR�;�-�.CR]���1Ҝ��Z�R��Z�(�a�A'��)�M�GB�#�f=T4� A���+V�LWğT`�k̽�f�	��єF��?i�$>�l��Cͷ��W��lA�_2oIH��_D����PG�A���������D���g0������ٕ�V���sަ<. xC���1����cd<E�z鶳PA&�i.��d\YM���*NAF~�	@RPC��#hH��7,�۱zO2�z'>��Mh�&P������<V��>�u�Ј�]m�לO'S<��_	��TI�|v*�b��P	������/bNb�d�[�6e���=���^�_Q��]�l�V;F��V�Έ)�)�W$�����U����,��M�c��E��~�=Z��rsX�<aa ��2%sٰ=�J�w��8H�l@�LĹ�63
Fxx��E3��t�T��[�$��/��W�3�G1���� u�8���
ƶ��ro���ŔTz��U�1�tͲ5<h6-8�Ps�C���jlxm^4�y���rDl����M3ù|�i����%&�i���~ #w��/�h[��H�*��m�C�������<���y��{���)�Ë��L��x;"���垏Ü��[#;a����Z�m�P�KOy^2��`i�u��g�#�ق�G�����%j"��պ^
�j�-3i�rPm{hT�b-��E)�]sn��J�Ӿ��q��
Ar�?��i^�O�j����?�P� �r�b�{�Yb!^���S}�c��+ޝa+���1 Q��������A# �If�,4n�on0�d"��X��wC?�`�W�x,��̅��]�O���Q��Dvl� xN�[]��NP~$���{[��4u�2x���D���?h�O����?��t��O�0�ȿABL����@$lQ�k>:�ioHvd��_��a
��#��)��v���D�ܣ-)KV�7h:�
�RJ����h���R-s
���c�~��@̡�`H�A����)��\������uʌM�`榷Sj��J�5���2Ń��O�\�p�(���'���{�� �*T�+'�����I����MN+ʲB�l/�99��P�pT���C��`�P~����ئb����⇶�
�N\%,X���CXR�|���J�
4�u�w��=6_��+3����)��������������������Z\�V:��dḞc�)����\�f\ph_!���8�[T��_?�֏FD:{[��V�^�G|�'��l6���#����p]�Z�O#���ɻ�ݼ�3�q��
gܕ1sQf�=ԙ�������=�r;��r�V��9��O+f��qN8o�����v]��]??B�¥��E���i��5`��+�9�ё܈P��T�����jA������|�s����{�	A�M����@za^#��HeY��Է�Zw�iw�Et��9E��KU7�K�
��SV��<�s�\��r�=�ޘ��[������f�k����,�[�wy����C��6�x�N�f<<��
�Qc8lD�����2L+�	�Ջ�t$�)�i*E��Fʫ��լv��%�<�c�G\��P�C*�QԲ������c$��[���g��\�0�zR0�e����e=V!>�	l��Z�9H��cm��kt��	���L�H׵̴�j�B��O��9vҧ��x��m
���N�����Z��wi��ݠOCH�\̘�J�%n��D���!:	�ܙA��@��r��+�N4!1��W�²�0a&_S� �וAe�Z����$��1rR�J�PY���2yL;d��ˈ��.���fh&�N �>'�5��"{����c�uB��4K�ыܠu5�$�c�]b{�)���Y���G��@yԮ��<t!ܲ�ɯ*VϤ��_���ȕ�B���E��Q��0-�"�K��D�����5�Q�_-�p9/	sB�����4���k%ƕ};~�q9xM�F�G�Z0��u�f��?4��Xa�����ڸc��#��jSW8O������	H͗�6�t|�ziڷ���1�?�*��G��a�;�$=�n.^CQ���\�)ӝ��n�u�NG�!*��0H�$�j��Y�p�i}�s�|[�}~&HA޴(W@����/���$e�z�)� �?,�<�/�� ��㸧Ջ♋�Ēwf,λ#���J*2�h��ɚ���/��+���&|�*�g:��ՊY��<l]�|�ͻ^�!d���Nt��^ )��j
W�����>�m��S�bø�Q@� �P�<���x|�K?�K����3f��*�_�uVn	pw����՝�_[Δm'ʋ�?;��Ususm"��J���6:~��&��b�&���e�X��������*S�][P|���}ְn��H'4P8�t�f��i�9~���:L��}��m*ULa��!�0S��|��O���$�C�:0޹�鳰�D+R@3�F��<�5
�Gr<��ܚL~�@�\^@��$�]�+�deR'�	5�����4W���q���,p;=;(��-j�����x�c���7��X�}IwV�v��B�N`4]��Z��J]�m���W��dΗ�a���0o�W'j�	_��M�ÞN;!�BF��0�'l����4����:�nλ����(�j�G��X.'&�ܖ�Fkz*���+E���=��]�&n�_��9�ٽ�� �p;����JQ�(��A�PN��ة�,�c�P5+ky���ų�d���D�̘������H�Ԭ:m�?i�I1��0��R�5	{��Ӫ �����:�a���e߳Ea�@OV-P�������7��S�6�o�*4F]��钼9&�e?��:v�@cogB"�M&V�*e�4���N��B<a��f�|?kq_E����Όm��r�9�F�Dە挺��(�W=(5�1�2X�.����)��Z?#R�i�X��;���>.�g� *���O��4�3�@�:_DL!h��B�w�0^?�BIk�Q$e�j�#��⋴D��i����4��x�k����3=;T�/-g���U-��p�A����ϼ�B�o�Y��t�����Ճf��{��
E<����0bq��va�������e���Rwc�K2J���|f��a>n���ҟ����CFQ�՚��)b}G��%�����OQ	���� Fs�&)j��0a�ݒ�e�V�dm�¹���v�X/9q�)�yX����Xm`\�a�,�I���Ta����!!����x�0��ʓH_G Wz+�w���"���Ͷ��l��9��N0�Yg�m��-<m�� ��'R�F�����̙����~\�O�e��'�ń�y��4��(�@z	M��mۦ_��~����<�r��z�[��z&������;��ZQc�2�&��
�PxN~M� ��5)�.��7�Ƌu��z�&Z�$y�.SI���j蠜�!^
!��%ۊ�*7�^��a���o#�+����K
�@�(�Q<��VӨ�3Dj;�[��MO�V�]X ��_�<~u�[9�O�Ӊ�"��G�ߧ��i�MK �{#	oJ���)�
%�����by��	��0���f��hGV���������(k.H(͖���\J~z�	a�Bl��8�i���x�K�]�f�Ej�&�E�Mo�[��K.2~P��BO�����w�mZ��u�	j�,�UX�Wg���-|�����"�23��փ�J����#����d��>��#G�{���̱�� �-Gr{��d�%��۳m���|�]Ì��i�Q���dv
�v�m����;v֪��y�G��,��ie�3i�=��v�'�%R*p��$��G5� �*T�9)"_oӒ-��S6��Pޟ:�f���?~�%H���$l��Fh�,q�B�o�m�"�/=� �*t8���}B�cQ����C��F�5Pqm��{3�1^��8!���~�%\֠�<�� H��q�k������P:��;k#6�4R`gF�(�=���B�Z^�0�U#�>���2���!��~!s�K�b���V��� /��by&��~�����_�i���8QJ�JͬO8��c$��P�u%���Z6	dd�I�c�2q���I�P�|!�ρ�d���m�ZD��s�~������59��S�SԮ[t(��\L��qJ)k�����b�����|^�vŞ�W��5��6���0��ͣ�xW�p��g�Д�
Ϛ�=�}����;�$�Ǳ�[�����N�S�gK��e/aq1�2�E���X�E��� U(������p�J)���X!��U8*��s���"��<�1�t�c�Q��Ҋxn=�SZ��[4L85嚓���ؠ�����0,l��еs�'�#I����Q���uF�%h���  ��d�n3�g���h@�&��#$��\�ʐI%Ж);�F���73<tܩzƍΑd0�}�͗�b���	�O$C+C+��f��ɡa�E_�br1 ii�"e~C��1�[�frԩ�PJ��	ȫ�0n�l �Ml�-$fh�Ro z�J�4S�� n�=s�>6H�9��I���d:I@� �N��O���rG�HMn<ζ`�R���`��X�k~�~�hA?��� c�3޻\y�p	e�����E��=5�J.l�M��E9�9�ܙ�(����m�sK��6,M���#�E�Lq�i���g�a�
,\ML���A�;��G>u�-�
7���Ɏِ���3' s�t�F{���M�wA��!Kw?n��2��;���@�':� �����w�[���w�)�Si���u�֚м�fڣ8��ၛ�В��ͩv[����-����5{�3�_���<H$��'^IO4�:U��-�=ʖ����vˌd��\'�ʩR��=�Q�b+)�g����IX��69D���N?B��p�vc+us����ι�A+��8�ʴ��T���%~�G���c�}[���:k�pe�T��]�~mn(�������_*ٰۉ��������������I����z]n���>d�1�'�C���ߣE���Դ��~Pˠ�9������z� lQ�RIȚ_��X��كuJ���w��9?��N��Z�i�6�8�r�>y?��"�&]�h����9�q�k��X�;�t����ı�Vj�hm��ݿf�Y�+�z&$�B:�cE�*��GdbQ�B�^����8n5x>�$}"֕�� L�x4t�o��K ����K�����?��S���qv5D���]�0�V�Imd�fd�AE%�n�FЉ߀�^W���:��"H1*L���yZ��?��uʈ�o�m0�j9J��ON|~쿭�H�Ee���l�3g���]C05ߴ_y�V�k�T(�ž����V%�I��[�9��M��5��ʙ*����x~�fR�Z^��2�Ӵ���Z)���&�~��C$W����H���;� �5�f��[�Jt
X�>������Z	,s!h
x,q��>�{/�/���8뿔�&�#����V�w������E�*$ش,?1^j���	�D�.�х�����182l@�(�v4�:.�d~�VH`)�G�y��.F��)�ΪE
�F"��3��Bk:����\�5�q��7��&%^�K�/���{��5
�.{�2h�;W�����,K/[�w�4x���f\ӽB���ˠ/��59�g�w��ɘv�����T<��W��Ac�i-)78�XzZǪK! =
�I��(��Z,Kڊ[Ne���2��ǽ�HWm/D�{�@���Ȭ*V+ǩ�?��+��"��f�>z�V^{���-mj9%�p�����
s��SԎQ"���9(��# �99]�� ���X�2������ޠ��Ƌ��q��;Jշ�?
>z#�`y��cT�\���<��sI4�����nr�@�(�ijq��$@���[�(KEA_�f��}-^Z(m��Snt)"]m������}�A"3ǪΆ�sg�����(�M���Np�cV��9}�eKn���/^�ajH@��|�AT�\7��$�DK���T6׫:�A�w�r�%Q��F��w|M/��	�E�\� db۽P��V�<��r���E�ٌZq*�ӲdB� ��U��������o{~N��W������"�/�v(������t������S���NQ)FY�&����pcip�/��"�Õ�/bj�eP�s�9���|d&lj�KB�a�E��J���ߐa���!$��@�����ftҘ��g^Y���\��tJ�&�ͭ�ɾbOHc4�ʐ�q�~)S��	���_��4�~@�@�Nk.BlJ���iFᎎ�Y�Q!4x����/,�9���=d�;mC��)\J�Z,��� �\܌Խ��?� -��E�����E�7��cFJw�Zd`,Y�o��5�۹4D�^v�$�F�FfF:癟j�a8;X��ְ�u���b�����.eE���c���1�M-�0P�r�j���.B�El����
��3�E:���]�E7�?N|���O4о���8�.��	O�  �>�5��F�E��}�Ko�5=,�4���]���l:�M$�r�1��x+�si��ˮ�����
��=k��i�+C�q�	IoE��dA�Ę�=��%�T:#}�0�@� �<�1-Rr��F]��Ղ���-b���dB=u�ж��*��F���"�$�Ly^�2�����[^vN]�c�5@6^d'����ȡ8�E�L�>��8��΋�">��'��u���wx�S"�b"�љA���7��YII~f�1�(U(\�"�k|>�O2�v�#@�����<����C�6q�6�F�;�i����!J�:����K����g��u� Q�����3ͱ#C ��A2��;�K�	#�M�V�!e���a��PI�����y��S ���@��|M��B�oK���g�D1��� ��.o�R�����]e0�L�1��ػ�0�q�����L��0%���pg��&�Д0���滅�?0U.-Rt`Ē<wTu�+}6��[켴<0-�]`_�֓	il~��}����xO�����C�O�����q$�h&�����V�=&��:�X+/p��w�}�)��k�LC����;����8-��_��
k:��^��+R75�I�/����C�|���߈MH�D�%ג�X�8�X1�f^��z}Cq�Ż ��bZ��g����̾�����ųV��R��	i�Ս��*{wA������S\��0 ��̧�>N��},F���W�^�I��4��jj< L %G.|�'�[qcD����K��x`�N�++�"h$c��&��My����>�'�I��8e�Y���q*����<��N��08_TwϥP7�H����솴W3��w�_��of���<����>] �n���H���;������S	������r�|h:�ñ��x����#��"~�$�ȶ 
���r�i��7miC��d�u�x���r�:�!��(�:�fb�<�N7Ax���`���]�Y�&j����x(4R���f �� ip2XgU[<h�U�䚼i�)�,�����v��*]s3�.�xP5�x���.���^����}���9�ug9�c1�v*]E�Ik����@��hs���yr��	��?h�5V��Xc�^��CL��9t�0\lL����`�;'��ܑd$��uwPђ%�x��»Y(��f!���Yα�?�+õ��-ME"{�v��#����.C\����ⵉ�5����I�.t烴L�o�q�tA-�阡Ǝ���6m0J���S�����cX�������2 ؕ�������X�����c*̧c���PYI{��EԂ�z	�A��cw�� +ȩ���a4��F�R�d�6[FT[k}��=ʽޗm�$� /z��N�͛�#�[�Ⱥ�q{s�os�-5�4?��d�$C\D����9t�˿���ج����c�>7��^�y3�����mJ�8K��Lq�	j�QJᨅ��p��ߠ�~���I0��VP��V��U�`��4�2���T��J�b�"�3:���~��$C�W�%�7
ve��j��L� �	5�[4 Wɮ,��QL��R�~�����_�p�)��Z�M�V]t��}��θ�Ғ�9c��� ��ݾ�iFx�*%V�7�939KS�m>M��-���j��^�P������f�<����bȗ����.��������u�s��77,!
>��.b嬑V[#ݔ��ϕ�`��=��Ny�:���
O�Ւ��8��V�\ �宯�=r>��V���"����vnbl����Q3*�ۈӊ�
�-N}�3r��C���sVwP���MxD(t��gh)kjc�ǚk�Ue&�����R�B��}��2�r�x�.?��(���<w���/�ѓ�����v.}Ǳ�����@x����yj!�mۚ6X��)����w���/�1ϏN�"�����2�u����E]˕Ľ���B�<�9p�y��������6�����u�`���H����7�|&�I��cKr�F�^3J6��=C̃�ԡ����l��F��C��=�b�\j鿍�]�� ��W혃�ƟG��F]o�y{$J��3����C��n[�� �D߂9U$ׁ�Ss����2'������zM�&������W�m<+xY.��5"�����y\:8%v��jA���J,ws�X���Ω(���;�2�di�͒�e������bH�Y���FZ!r՟x��hQ�~�|W��(�1;uj7�̩T�)�VM��������a����={ŝ��|�JU�G;��=�&ʄ��1L<�%^��4� ���H�A���N?\0�I5=6�`�ۇ�w��8�p���!$�l��?�t�հ���2�悟�˿s A�+V9c�G�C��C�_l#-�5�(;"�v^��[%��B���HrB�U��H�_�&�oNC�qґ����3�6��|� 
�J]\�o7膙GD[�nr��>{�CX[[Ut�A���[���4���n�mbRΩ�X143>:��y(��n�R�<x7��BkL�n�Dّ���l@n,�>�@��%�[r\��&R�OSC�N����v��?���#@�q���qI�U�+���}m88 Zؔ�>���K����%:7��G���8����j&��q0�-##v�{-�^S;�38����n3� ��l��$>��50��+b9p=6��%k���U��9s��7��:�7\Q��I�26�u���O̤}����<��>��f�9Xd����a�ۏ4	���D�,�a���W^��]����?e�������t��	�*/�	�����k�����S����LmSw��b�sFjkJT�`r�(Y+'Tf���9(����B�;��el10�=�D�LG�R�Y����P���g�����	�o�����H��c�l}`1 �7��6��c�= {0�꧌!��>3�`�d~%�Sd`�����qr�
�A�l/���f��������Tb��������V�܃*҃2�g���h<�ֶ(�Ui�� �̆Ǔ��q�<F�@��s��.�x���H<%��@#�7���U}���A�V�rMk&L)�XQ�U���w��w+�9D����/Ub�{ONo��:���ՅF52p��1�+"&�
i�!��8�� ^g�������:���15����Fa�AL���>��z��~�<]������<t{׀�u��,��F%��T ����)O]sS�aB�u5<�"uk�L�ks�P�ſ*���] �/�M�H�=���)s��9 W�@�)r�	}��o��Vj����ZYm����=\R����-�����M�1��lF�Cl5��UK�"�|/����,�-sV��;��s�R�.�q�a��5�L1�/c��Z�J��7^���=U�;�wK�m�b=9$@C6\��jh��d:���g�c�-{'���7��ڀr��}�,�(�k�"�p��׆�*��ɻ�"�Q���E7�Wl�y����q4]î�%A(�<�e��
��9�m�H�M��.�4�����u�(Kn�Ԋ 1$��)�(��$P��,NUϱ�w���TE�'�[����wV��P�g�?�iB�µ�I�e<�Z*�����!� !��θ�_���5����_������A��&��9,�U���R��W
���)�[�����ẅ́��J�I�٥�L�, ���A� b����c�8ĴE3�h̩bz�f_���:�tʔe0m��qQ���LЈ���Ƚ���^+C���q��U&滸�q����T�T!��7I?���3�w�����Cд
6���s��ѥ\�I#�u��i[��Д�D0�S�p������s����4ߚXG�$�����4���z�n�1'��s._	��s���r���mIW	G��T�������O�:�w'�> C�9�%wX!I��WD2��sV�x�w�.蓡��J�bc�9='N�]�`e��3�Э'y��5�T<�ٷx�~>V�d��X�0u�
z��!��'ǅ/��"K!�-�5xz��V�#��Bɖ�a�����e�D31�C�RU��:�G9�#N�Օ��\��r�a��\b�6Y�w~ݓv�R�7����T���D��b���ݿ q�^�3�!ҙ�~��}������(QH� �V�#p%�kn��7��p!�װB��e�{��8FLz�ӗ�`4��4^�[��$���Ure�J�|��݊�?x�7Uܨ�˟���+���'T@6 �I��nf��j1�c�67<3�$E�������N��f$��?�H����Jϻ����.cѲe�Gf��R{.�W]�E�G�u!��s�"x�rg�u]�"��w���� K�F���4H�
ųfƿ�ɹ_\Ӱ;yq�� �fP,�L�&-�;c
vp�p��P2���u�~W!�xݫNv2k��.8��J��L���D���Kn=B)s������B|4 wI(�`� ��ח�t��'�Q���,�B�x�^�~(���@h>z;ȝe�71��z���Ǥ��e��^��=.b������c���ׁe2ZГM�X)�M�J�Tg�6�-���=s��.���%��E�������l��?�J��=������1��J��;�&�n���nV��*�Qy���jI��x��c$cB��������0���[��^[9��AZ�q�1�F������q��՘�m�~�
Ź��v]�Ď�t�į�:X������׬5D��G��IH��N���^����t
��W[�۰{��j4?}GE���ؼ�̝��X���m�?cp�ٿ��V���|/p�A�9�ʝ�vuө��j`�B-������@�J�7nE���lg�n�	`vs.A�7��p��?VfL�{a��������.���U�9[���!t�OE�'=�%��풖�Tx�S�qt�����Q�f=`E�M8�޻���B0�ƕ�׌�z��
=��ud��ZJ��6�W*�?9�!��Xw�Qk� �jW��ڊ}5T�(l�o�j�ײQ)��=�/���9��=l3t��ŭ��#�]��m�s*�
��3,�.��b�����(봦\�L��"Q ��Ͱ^^��\}�!|�1TQ����7R���hNf��w�6�Iy�.D1s}Z���v��nךw���GѲ��e���D(�2<t-����76�;؆�p�qg�G���?ӟvٔ�:nO�B���P�J�>ֻMP�e�췣�yآ�a5�伜2�Ro�� �=��F�r�g�t���b(����+?��&�C�p�,ɹ�|�@d�.]��ti��ףH��o� ��Ͷ?{ӂ,���e��a���b��i�ɖ�{���ET�������1F�q�p��
�vP%����`3w@[ēPr�Cfj?�aJp ]�$�"a5���Mh������X~���.��p���@~��{y3�I��C0��*�2�T�=��'��уH���r�)�8�5)�w�ʯCB9�`H1�c�'/�tH��
�n�B�9���x�c���'��癩1��C�g��w��e_�A7R��XQ�EuSb�n8Z�c��������O��ժ�8�VqLl��?�{�->� ���2Xe�@������c<���������ؓ�CZ-��/�a�Y	� (�ܡ�
�j[+�"����I{f7�q�X���)�,���`#�9��O��<9��/a���`H2x̕M�UK��7�T^�;'$y]^a�7ڟ�Y!bйʦ\fG���C��s ���h����$Br�X�i8�f�n|�{R[;�g<�q��݉�N���K̼��Za����NH4u�l��	�X���~T!��������z��t����q��$:t���7������A����?,���W�V�4h�D���(T*���>x&�|�����\����4|�](Ib�el)q9�&+�-�g���#��2���c��p1�^��* �w.��=�eNEI�c���,�(⃋�\�����b�w���EN��K>�8�E'�ev�%�����֔�������V�q�f埢Q銔s�xv�Ck��nlg���h^Tƪ�j�A#ː�}'՘Us$_�YjZjUgpj��K'�-� uR����'�^-D{߿���$���?�v��n��Qb1Y
��b��Z�A����چ@c"/�0���А�� �QF�i^��lav<� ݂\ҖW��ueM�܂�v��0Vٻ��b2�b��S*�Uy��xC&�_܏�f�W�us�G	�0aoи;	���BΘ]�5��(��NFyb'��b�I̡|c"�9o^0'��6�=�2�Q�q�,��s+�D狎�؀hf�������(x�c����xb�u�YЏ�M�?쟰�d��~�(:�,��t.dxF��1�P�"�B= ��gj���f��vqI�kb�<`婑�'@�3�rX\�r��*�RH��"W�͗އp��.v�+?��mPC�#������a�B9���~$c�)�OXR�`�c�����+�Ui宗� ��@5���Hw���K�7���cIg/��������y�������1��j�WPQ��7��^o�trA�g:�<����O�#����(9���װ��PEDU��OC}�r�2CI�kT�V�#���FwCK�3Kp>opT(�9{��K<g�)��Ǐ�au��e**�x�g�R�7OF�z̜�ZA�N�N�?u)�(����j%��p}�I���0�+�����9�ɵa��jȚ��S��W��54��\�꘏+�����d��K*fYJ�p�w��~0Fc��;�&d-ՆMx++�"�hӼ�e�j�xG�{�F�zi�$�g������B튧�RQg�=�`T��#�4w�^ת#Ti��h	�e����z��T�P�U���\��&� �`n���:�OQU��Ĕ�P%��o���9xzɢ�Q�J��~�Y�"���V�W�}N�3^9�Ty�B�l��ٜ�%5I��\m�pWnfu��l�~�K8���5X����t#�唸Lh�����r�o��_5�����ݐ" �����!Җ�m�"i�Q��b��d���$��~��y";��ND�m��J����)2N�>�E��<�;�"ެ�E��ATvy㒎	鼍ce�:���7�Rr�V���P����$|j�5��Ҏ���˝�iS1��7HPx�'�g��S)���]_�Q��M[V�25�V��cqm:7����¨%�
o�4��A��3�rƕ.�T�X��p�c��
>8�b���N�
���9�i�a�R`P:�8��2fd�sx��5�og���s$�ob*C")q#=j��4����Ĕ�"T�oZ���U�>>�����ѳ�(5���t���4��t^�ݞ2F#�(��m�6]2����U��rԨ�4�����n臃�t$�E��U3����jn/�3�����p��U-�Q'�t4޹6�6?��*�8_9x����s)�DxL��JGG;�$Vv�rHSR@U�Ƭ5�RJ{K`!x �[��$j�D����tCN܍�96��gY��|@�(�K}��
Av'�q#�c.\aCySi��1����BR��>�:8UN�D�w^�]�ͧ%Ԑ��f+=}�~>uM��_�7�E�=���(H�J���ɂ.q�ۋ?�$�����n1�_��w���o�v�j����ņ��Z���WeU �CV�?���.~�Xo�_��a�%?��O�����U�b�Wd7Ֆ�L�.K@�
a Ǌ@,s�3�5}��&�k�&���P�����w�,߱�KM��5�u�ń��-s�9O�+)��2a�'G�I�ѮEG�."++H����-F/�j��A	̯:(�M��5�J�@_�B5mI}�?;��}��a���|g��fS�M�d:�|�����ASŮ&����H�}�P�&5@���hHJ�;��\զLG ɇ�G�~i��d���cbo�Lkhko�����C��)EΙ���L�
�"�v��z�-O5M�ͻ�묣WR��z6����|Ϲ�>|����|n��,:�tNZm�so	Co!&��b��j$��H��-�Ȱ�'̛�,�&-s��K���*��ΟI�b�'�ߊ�i,�f�Ƥ�H8]�	^N�f��[ |���$��c�>��8��Y���4�?p`?��g/p.d[���9*���~��*��
֓نʺ��Y�c	 lnp�#J2	>� U���jq�/��M}��pRB���M���=Ĉ�u�����kT�ZD�\���:��h�j:^(���C<!�9tqP	;��:"E�����&��A�i$}ɕ��:�ػB�� ,��7����2����-E�Xr�Rf���s ���F�d��Ɣ����������˓�\����ka&�68�Q^��p3������-9������5`Z������ �K�f�WsX��oHQ�Z��˟�.��V��S,�0�ڠ/��S�ħ�㈆�*Ex+7���G����&ZG�&��4rԫ���C�p7�t��9u��넳u��#5�����������;�`��&�h�uH%fc����3~G�:�C9l��T�>�R�V��O�%��~���n�~/��j�O` ��Ǭ(zP{�U�4��ߖ��w�t�߼j�K�jXa���@u���+B�G�r�ti�q<�/� �Wp��J:���W�Rgq�:�2P_�'ir�,�
��4K�;�1|�CQ�j��7H�������i ��E?𓤿_�/5hc��6�����ޤ���-��)`�SуV懊�
|&;�V����#�f�W����43{�s�|<�6 #�
K
�oL�x~��s�}����/������#�n#w:����]�*3�ö%�������0�&��3��\���A[`� UsX���$uA�h`8\�BF� L띶w�x�SB�E�)�8�i�3��#�[᪏��7>��Y���R��I�KbO	��e�E	�[���7��ӥF�� ���ꝒǤ�� ��kH,�%l,cT�d|�G��� 	e���QPWճ�ۦ������r�NV��K\a�y��n�}��j��Q�*��!�<�����/ �0M.�,����$�d��#��
����q�`��E9�O��(�R�?�DG����{����BjZ�i�l:�,�+8�|T~��g�{7��\��v� bL�F]�%%A�S8�u�w�Pk����#œWj�u1�<1v����hCCIFrXS!F�����4v�������=�c�+~��,��I�����\�F���j$�0��Q64�_6Y��w������@��h���o^4�|�+-z�<�<41�H��C�m��� Q�������{O;���i��Vۅ9��Ф��)��'�����M��Z�2G6�t��90����lQʌ�J�6G��	>�en��T/S�x��tB�f=u�n�L5��l#u���.�[;���}�?����k2w��% �&-R:V6��Q8�,ܣ�H����[��Ȳ�Nw�vA��
��+�]
�FgƋ0#m��8:Lf� ���m��H8��������D\k��ԍt�Z�ܾB���H�m˲�2������ҊA�Փαҫ��-�(��f-{KnZ�.�]��;j#M�rUOKj�e�Y�Qf��;�o���"~{����H��_��o��A,�x��Z	�V�}	b������Q�"��	��}ɏ���x�]��Pᗯ\�#l[�+���ȭg�+b�Y�T嶔����H��U�<p��EЩ8Њ�"к,;�`*�:�H�W��-�����e&z]�C3e�	�=g��d�E|QT�~0��NN)CAYHK�5�f��<�E��9~Kмj�Z��iyhI��g�{*�}��=%�Cz����B	�}��J��T�R�i�=z�[�J�O�Cf�"؝ڄ�[ͦ�������DJ��Oı���h{M�p&��I>rN��=L��ߝRm�����۬[�=�ǎ	�g�}��\�P��(��Db��,��iS=y���`��������}�^�8�Q��	E1�<�C�	"_kz`G��ng:�<7ö�3�HM̿ڐ��L���+(j%�^^BO��94���8��QE�����l��~+���{¢��GC��P���թ�f�a�92nT=q���"���2�j�F\�IHA�a(��C���X�u4�ܓ� �{��6�S�8�KA����HȐr�.��}��dG� aF��)�2��=T�|���n��|f(:D��Ь	Q=X�b��KJ���T1,������d2߫�\8����> o3�Z|��/A�af*c_�#\'?�x�)od켈��u{|ך�[�3�B�� �����hZ �_*##�0���YQ6[S�|�3�2��G����� m�Q�Nb�:�p�0H�.R׵_>����X~���&k��{�&�j��
(���!lY;�qu^AD5�Wgb�ڿ�d��Ԩ��%}z*�O5�ʕ� vD���I4l�ww÷w+��!�jS`&u,A����FdVu'<'���������H'�
�^��,r��@4���ڃ9`���^���݂+��ex���e��A����m����1�o��C/|�l >E�g3d_�&�-d��8i��&�z��^m�����U���j5)�����p�e1�Q�?���.���"9���\���Ϸ/A�rC��L�&��+�����_���Ƨz�&���3%��xć�M���s=Kb���*0m0_�ǰ�O�<i&��&�U�)춒�9��*�,�r�BFc�6k�Ø��m�\��������%)���k��i��X�21�3�R�b��h�"�@'��}^��jX���[HBW���:�z��q$��z�a���>+6a��I��%ʧ�u��>d��+���sŤw�\���q�V\'�'����0����Ze0�=��K�bQ��+��i5��!9p���-�.W��뻅N�3*{')��~������C��;�������t�nQ����� ��LvBR͞C�C�7i�e	��wi�f�a?9&�OQ�ex�
pq�$�y�DWe�ڝ��s��y�L���.��8�B|~�����o(�8=Ea����������ve���H�D���g�����r����B���P+^"\�%�}��O��c�9Ǡ��G`:$
�h�V���GTocb:����kM� C�è=�z�����A�?)�o���DT�������v��%����ǂ�2�b���0 J�a��>N�$�������5G��X���9lP�ʉN���ꠅ�����ۑ�������v�����z���lzo��������Lٕ�O�e��r��� ]�U���Ne�֐�yԤB�y����j�.�)�<U��`����9��>Ww�O�=��i�� B�!�{�}�%�w���]�3 ����G��Bhٯ���AA*�c��4��8�Fp̹�;�¥b���1+[�)'���^d�IXH9�r���B���vR����	˃#A���F!y� 
br�j�մI��_� �O���J��6P��0��^H��f��
2�B�T�N5�˙ a��x���F�kU~s^k�Dq��L�M��b"���U�gs�Ìa0"7ӾydǢw�VBCFa���]���L)� ���w#���R�U�)�µϕ��Y9`��b�c���j�7#���ҩ�)\��J�r�*q
s?*��:�s	�O�;�\�x�?��� lx@�\�]b]?��ت�w�)\@�����U��-?B;Ys0�j�+�3gX*�?��������O~m���Vֺ�%ڳy�>����[D̀�5a4�3��O�-����;چ���J�V_3z5������H�J�j���Xٔ�=Rz�5�S�p,y��|z�ig�-k�8i���v��u�@tg���I��(�O�WZ�f��=��5��%��Üm�7�<nq�E���H_H9G�z7�1�`�P�>��K)�_�]��H�J��̩���\Scq,.��b��d�r�+#�Di�������MrHH��6�_f��I������}��P����J�$�����	
��"������;!��lk��N�1\�C�H��QLvV�"I�o���&|h���>�Lgk����/���$`�M!Ա
�Mp��ۺ[�)�YץT����δ8±G�Ɵ^"�K���z��V
$ۯ/�QSK�84*D��\�1�#�Ƀ���D��!�� � e����Nj1�<�j������O�G��j� �m	��ď�w�E;BE\�N$��4_�qB/����vDQ��?�ѭ~�4*h��G���rbI�PuHݓ1h�*���k��L/*���m17�k�9l�%-VW���`/ǁ���з�>�h�$ⵛd���,� *�j�B�t�C��+�k���)x啸��$�I���m�W�	l�ܧu�I�Yo#ph�=�Lth$Y7R�k�z���$"�J|�%r�A~V�΄��v��,���K.�5�ōw�F���3��?����¼wp�!�!?��ID�W2/4����>�o�w��tvM91�E�ULo�0i�^��|𔓢k�����PL����G�:�!��O�"�8�ܖN&�(�zɒ!�HXzs��?I&�!��mM���8�07���3Q�4;?h��6���s��Ю��H0;cObM|(w��-zx+@���Q��3��0T�6����y4�v��a���z!]��՗͎���,+r�G+f�"���Q�b�q<��[s���w�95K��gMf1�H+����)�P��*f��7�W��� �p]��)z(x?��e9{�p���yA����+��T�>�׫7Sv���V~d#��H˚������?%��S�b��g�|�vW��2��3���RNI��	�U�H�zǺBJ���҂q��%��5�ߗt�o�<�t1��a<�"��~�]�o�DV���GǦ7fu"���C�5X]T4��m=�j~�yn�rI&{3Z��m+� \/ו����%�vC�0r����DVz�b�.Z\7��l�21¯�kw�l�S�c6�43e��''i�a����k��(�/?<h3�L+)ٱ��o
Ï�T.��F���2��
w�8sA}� �Q��Ӝ��Wd�mj���E��;��@�|��8e4�H����q��,���|�w�Qz��E��.�d�n����6Z�>,W��b�!]�!-@��Q@�Yep���q��?����MЄ�*���ʙ�U�6G�%����u�O���FҢ��ޖ�4��8�f��A���8�M�Kٌf�oݜ~��h���\�*r��|R�<ӏˠE�H��y)DB{H���:�ӛ�����q��Dj�Zq��	�f
,�O�B/.����&g¡���7���Y>I�2�`��F��bR�wJy��Q���L�hH$C�$��������eX-K�:ip��$+�U�竾K��&)C-s�4�<�O%��;E���h&�[GV~(�ܑu���C��Xp���J�#������|"f�5�D��F�U����r��=f�_
�j�~�Le�˄̷=Qe�r���K����7�i�]b��%�7��I�*���G���C�t_����=��3�2�?��ի^�Dv�Ҩ�S���9gɩl���τy�L�~���߀%߅��[�@�9�<�'M6��φ��x��7��.���L���,��^U��?a�9�9�s��6щ�Ǯ��ua`I�z��Q��{y+4�;��5U�g��ɤ���jZ�h)BU�
F�n�������R���^���� tb��,��;�$B���T�es:��
tj��>��n�He[GS�tY��-|flc�=���z����,C��8j�5N�N���&�:�b^�^o��;��pz3��%�U:n�,�R���zl�Ŗ��TB��)�K��g�EY�O�(A��ﲶu���]��#����X�b�z��l�������dO�,C���`]KJ(]�֞��8YqV�M�T� e�HD&B~�~^�(�Q�vaCFB���GE��$tBHP/��D��S�l�vfˣjr0J[x��Г�5&�^�P���ϱ�����a�VK�^���)<((Tk��˕N���X��8���J|��rz����x�������7�㕨�%��	=��M��c�1ø�r�b>�O�Z�#�K��ѐ�X	Q9�i �&e+�����f���WƾOΐ��!ӯ�ᡚ���YH/�V^�e_�C"�/���J��M��Вt�s@��(m|R����AL7���YA�Ϧ���-���qK-�/�^��l{�[3o�	^�/R���ک2@<��|,��,�Pe���up1/;�I�ǰ[s?2��D�;$!�l��D<%��"��g,a��X�Y�Ӫ����%����.D`v�m�r�i������>:�B�Ο�4/�^-���ŭn�o}�(1s�._[W*��nl*)Hol��%j���eӶ���������YA��p&F���o8���C"ج.Ȱ��B�{��O��n�y�F���Aʀ��Q6H�!�[Y��� 8�C��n�xQ5��&q��d��%�2�QM �%��⨤4\�$��>�4���Ώ[��Baj�O�z����F��5�ӚO�̽���l�o��R��� ����'���u�|��rM~�A$�2?T_In��\fH����p�$%�U-Z�����ħ�������w��V���2b;W\WsA�T�ds*h+'U���h_��U��9D��PҗG�k9�ۉԵk�z�6�?A��R�w�Gif�z�	o�f�ؒ�Q�1��Ϧ��Ђ�?��}�m3 ��v�%+K/��=�,������[;RQp��BN6��ġ�O)��k�Bjܵ����	�����f�~���Q�*mf�@N���]a	�a�s%�z���:�MqNə�z^��h3k��m�;�3F/^�F��	E�½>נ}�xpI�t�q�-D��hv�_g���N��|q�E�D�|���i� _�-�.b��r�U�M��
�r�A"�f��HЉ�+��0�0�ew��ذ]%t�[�t?�jR��Ӟ2!�ѵE%hB�� �M�b�J�VsNK�8�v9���;V�R\��m	%/�z>��"%x��f���iSB�
�nH�#�-�E���=R~WS�P D�)i�&R��m��/zݵu.��a�j���.�8����&�C�Q~�`������

��aш���E�R$�f2�o��#�G볪��+VOh��Gb�ήS��Z��,���؋k�Y#� :����A��%*�R$w ya4�{(�9	�!޷����XtL��LN���i[R�ŝ�Ho1j��¤��d����w��~ �3;A6��K����Z���Y�X5Q�%�����'��!�Ij^���>�>^���1e)%-k�, 9K"{]��0�.X�
J9�QD ���O�$��y
�g��8�������v�5GJ�����A�g��ȗF&GMt@��[��@��:����GB �J�}&�~d�|�yz�^�M^��5/)ǌ[hE�٭�������P��NQYY?������Đ�Ԉ��J��*�#\�8�!3g���	�����-PE�KD��(X��D�&`����,:�G��[E�5^�ֹ�>�q��`'��B��Yj�C>����`�
��mꮉP����Т����{�r����>�Ÿd�,�����,4�_��]֪0a�LC?&rI��x���3[EvM�@�hs�ׁ�5�4����2�m�0I��}��}K�1|zej�p�=)l� ���D�zҾq���9뤕b��W�܂���`����l����tiVc�V��	fd`��AHo0/D�?�.��4�&hCJF�sB�/��p
l�:�O-�8��$;�s)J��+��	�I'&�M���cZG��t��S\J�Y"Q���V*<��R�ɰ�i ���R9k������N�5�x�2��(��8(��qw�B�9�vH��c�&Й>|N��>|�H�([B�\2C��JZ �Kȗ����-�������Y� ���#�Kj9����B�LBQ���֍�puT�x�@Tn�kj����!�#.��� Fb���W<�VRD�돹'7+Wi�� ��;�"�i�5܎vF>�y�h�o"Qy_��C��|�Z0��T���3o�>�E�+R�,&ّ�d�8��)K�H������
1ꀳ�W��9��.���n;�n�%����=�Ϗ���a��G��m}3w��+t��#sY���4gA�ƕ�Zb�P�����
)3�ӓ�������+���vh:�s���30�=��ֶ�/�c�oi����������[�FA�=NtJ�����O����/6�q������b�/��;/�Ad�vg��Y��05H*C�D]�f�szȖ��*Oc�L��9�n��IԲ�#>���m(6��Q�SoU/���.�)Hku���J>��Mg�E�4��ʧꄍov�l��F{R�4ԟ���?��i��I��'��vR�q�C���V��3%�`�"�A��N�D�sv4J�8cel��vſ�v��};P��/W$q�#�a���,�E���k�H]���<8�c�/i�p<�tAt�:s�ů<'�s�L�u<�Uqa��>v��v��3��K,L�~_�	����1�'��I�c������!y$s��F�^&I��/-�9�8�it�>z����G?�F���*M�4��}v6^�+���a������`�r�7/�R�EW�Z���:|�� �BM~*��6��lMKø��(�F�����(l���8 �z�j6X�0B���}��á�k������������p*�O?%�x����ᚱR�1 �-����<M[��?Qi1���O�T���qD8\�5%=��F���HcGF���c~j,�z�k�p��o�q����X�ԫS��Ⱳ4���.���uZC��hzz�p��ﶽ���e��D�c%i� �۾��W��?7KKݭ��vjM���t�Aށe��p_�d�d-`� \��k~n_=m��G�E�����sX�&纻�<j�*�hD���b<I(����$ةN�8s�Q4��i��MA)1�Fo���D�=/XeW䞕#%]�>K9�3~��p��P�F��3HZ�o鴾��{%�p\�������^��thF�lc�;$��g`����N�Z���0���n:�n@;�T��\�	���*��y���z'�u��4�'� �_J /�*��DպZ�k����9nֹ��D�Pm���q�A=�3����(�ɚ|�.d�s��9��Y=�P�,��>�2W��y�@��=��I:�O�ڈ��~�@tC"F7T�r'N���k����.7���ύa��2�q�O�[�a�i��Ld��[��m$��f���llV/����A��S�v�;��了�ݤO �5�j�:� 0`���^
-�u(/�6�j�1���r��P��&��L¢�b3�*��g*����e����&���� ��H1��M�|���n��X��a/�@�v�W84I��BM��N�̴���U��D��L'�ό
_I�5G������ͅ��h?U�/�W;��\rlc���ȑ}�j4#HA��Yr`�ն,r�D��'���1����ۃ�9#a�'_D�`[v�+�/k��G�A�+QB�/��5\hxrzQFEHk�pYk�
=M�j,ɜ�R��:�m�O���^�mg}Xu��J���Q�{�����;v��PEԪ2c����X�s[��Rg
5�������8��ntI���`�?'p�(} ���Q������Ch�h뷿>��*�VD'm�A��0����RYP9�M��Č�dI�Ooh�Q�0nH);j�򄱼�B��!h0S zR��  �6>�-�>�88�_��}��A��m~��Y��3�����?���9N��x�K��10C�=�`=Y�a��$iМ��Z��')t��%��.��Ms���,L|]���~ʏ�jG�7 :��*37�T/l8e��k��!y��1��\�%%$qZ�0��L�݌3�����W�qbL�E��ק��n6�.!%����I�ϖpp
�i�@�v�N���s�u���e>_��[ffe0A��Y.	��Z�fS5�_��.h��������4����y8�P�(b싴�R�6�7�Na���ll.��c�h{��U[�"��>�'nh�ih"�����ྖ�7����T�_�������q�Pp��o����h
��{)�w�8��ׅ�t�'t�Uڗ�24Io�)���cѽ�>�b��@T����@�#����-�&�:e�?U���e]Ob����>���h��9Ǟnbդlno�H�x^Y��t��-ItYK�#�:�mߺb��H�	r��^�F��Jd��ʔF'�fJ�_/;�k>���N��+�G�����9�Zã��w�
�#EH�z]ǲ�spw%�LGm��ҏXf3Ӫ{�����t$Tz�w�&�	�����kEɆ�~'�����{��6��SGj��)��6a���wB�q���<(#VM�����Q�Л�M�iQ�z1��J�#f�1t���l��+�Ư�9N��o�����b�쵂&�>M���KR�K�H�s
�jd. o��U��X�s�z'_�&UPwLf_b`B�k�(���N�_��#�Y�qZ�jOt���ٚ�f��X��n�θ~�j^�
Fv�X@��,t��w�5�p�%�W��O�U��=N(��^�F	2RY���N�I��X�(k��Ҟ�Ι��e�Z��u��@�5*�.">L�P��ב�/���[�gk�􃖮�"#dT�]<ox�B�_�PL�X�[Na��W#���v��Z������F�z@�Ფoy�UF�((�{��RO�H�f,&������N�>e->*,?V���P����YOa�zAPQ�i��N��&́��<�Pn�}R�nq�ѯ����6
Kft�]kD��l���V4ґ�9y8�`.�H�\���C8��Kvl�}��k�i�B*�[���ӷ2�zO�w<9_D�M�E��}I�UcN�_��E:i�@V��r���K�5$�d���Dl�wE����.v��yL�����0U�I/��1~ۉ��g陳}�>�����O�O�����I���,:���ةbr t:�38\}p臭a&o$��֦���1&#��Op�Ш�<[�ě���k����0��LC�����j|��^��YO���ϔCw"�[�5I{���\�{{XSA?�Jc�Ғ�������G#��]~��r���:�O2���bjO��s��Rs�#�T7�@�T@���u�!Ō2��ѻ)O�E�E�$�8�[�^а��������F"�q�2;ݲk�Nf-����	j��Ȇ	1�]y~5���+g�s_& Ҍ����`��8��?�y�j}/[�m^q-U����r͖�?$l�TE�nӂ��^�Π'^Z��q܁�5}�Do3pv|���%	����q���@>����5����U:8Æ�ϔ�$=��X�0��������۪6�A-��=yuL	����2��G_�:��L���.���n7�9�j@��r���B�#!q���N`��3G�l���ڗ��;?�1#E앴�;eӪ��'d��ᬉY����� �f��x���0��R���8�@r>+��2U�ƫ5�	��:��_��+\2���S"�ȍ�W@�	!E�y]��O�B$u��8C�DI�S��}YS�)��q�$(���]�k�+�N>o��4c{4ɛ ���.g������]���I	�ӇU�`K�z���}0�B��U�H��e$��N{�L��@]��c�ޣ[5BX��G}��Zg��-ˮ�* �����}#�u�n��E+�G� ����U&��0A�ĈS�@ .7�y�
���Ai+wD����_����[)/�"�lA!5��ǿ��7��)nl9�P�0C���{�d<���������.lPFr�3N8Lڊ�.��0���]î��Gh���NB-��q|*7�Ub�W�V|���̫�^�x��x��> �Aj��`7�
�zхs# ��*�1��+�ʑ7��u�|#�B�(���ş�u'�4Ҹ�M�;�	��Yja�S�2~U1j	�
�]q�l(7�\�gӬo�|�T����c-�os�<#b��_�U��m��=�u=�s����ݾ��F���ϙ��a���_9��mc�>w�]��F�?���b_o��w��hN~/:mo����gF�J�p�#-���ң��,��l�v*�PGi�9�����q���}�<+��S�C�R�^<R��ng9�ܤ��)zmz� �,��^Ƥ�t��U4�|e��2�Z��
~��G�k�+�`ș�wW.f�*G�$#>!L'��(l�5�)�q+��]��%]�D��M��.W��3��--�T�ɦVP�me���
zd��8���kkʌ�e��[1�������<�'��ErL|��*��5������i�'m�"�H@3���c�����D9�\�o����W�k�78	(� ��_�ؕ���Qܥ����M�[��z��>���Y�`߳Θ@�72u=sL�8���CPO���Ws˝�yp�NrX��]�ff_���B�r�L��N��P"��y�f�$��������5Xt�`��`Y�����b�UKs���מ����N�����fN��{�s���P�2�Վ��v�s ��np��b�X�߹��#�Mj��S�M���,���J�M��Ff��Kfjr�N׎}���6�G�([���Wr#LUSu���ɣ�.�0c��
QE��ۏ.�F�Y~���*��A�׻�C0�tC "o�nO�{bq[em폻�jl�=�>��@�I@n&' ��nW�tfAkr�����7�%�;�%=m�dT�u��Zk�Pn#J`��dwԱ~֍I���#??����q����pK9N�~NY�?�0No�}nװ��,'#x�𸣴;G"@)�R/0�w��G�j��4�׋F���<|ن����
g2���붟�O9<�i�*�1[���*�4�5�ռ��7���C닀��91ՙܿ���/Y�\b��%X�֠������P,�q�$�mu�Z�zfW۴�7	�������3̄�6N��+r*�[U����o�*��Z�O0��/����mj�H޾]
���z]h4
徍��e�b�E����G2[�ĕDQ�����pZ�hʏ�ƶy]��0��y�k�Kb` �'u�-O��	!C��?�O�v&Ջ����Ħ.Q�[7�IP�`[Ld������;������gv<�#��#���G��̲0����.n�~=�K�-5kwG����m��VY��L[A�n�_7�'���_��[��\�e�3��q�S��
0��R���CO�#�x(��@�½��lƷT��g"Ƥ��a���>��cX��$�a��6g&b�M����u}�$V�Z���%G�aA��cӤ�,� ؏Uv�ve�Zd�ݞS�l�YP.�%u0�2�7�
���Ytz)[�q�W�)�.8��Z�48�L�\���6}z�X�	y�� �qI�A�5ii8�Ƣ�U怺�%[�wl�;̳���oZ&9��l�=��;��iA�O��s���=xA��T�Mv}'��?HW��\�(=r��v�p��6�3�We��美��щQ�"(oe$��L���%��w �8f�J��ލ��]. d��4�'��
����C[� �#lQ��*�1u�+�˰ۆs7*�`Q0��];ۜ�/�:O�D�����������3{@��@���Gs�e�\����8����
o/o(:Y-���~�i� Jң�S"����!�?���{ ���×j�8�p7��}ܗ��{�d�gۏ��w�yV�> *��Q���ce?<�5,�?�>E8�@2����70(������?*��qL0d�s�$;��M|���v}9E���~���JG0�C��8�@g�m慷��1U�!/�.d 5�X��4qi��eH�3��A���/[�E�dAp�|A���RQI/��~�[ָ����S�c�v��g�r�S�Jk�K����V{�_�S��)��f^�G�fCa(�wlW�k^a4u%KE��`��u2ë����]:{����S���+�b�Odl�8�6b�v���Iq"��d����O�G�U�� �'b��{(�)��2�9Κi:�"*��S4����2����3W6Ur���LS`���DҬ����.��^�ɱ%g�x�ڙ�]�h��Py|<�=+nh�> 9�n�st���[�jyGݒw����i���$�wp ���;�$A% ����l��`�4XEH�I$u�C��&4�܌��~����l���`���Q��{"�K���ܚWX��ym�4��N��ZmK>ȥ)�1*fǭ�LGd�ȫ3R��ohO�;�7X��BTǎ��L3)|�������`�I�~���a����l)F��O����C����ٳ��4ip���g �\wŚ��#�Ym��=t�u�V��6�#������	BՄj7����[��H$x����4����Ű��b�X�׬|���A��(.-����f4 ����2���wuB	0 �ic쥖��BG����S-���v�l��e_bp�F�����~Qa_���S���/:Z�k����>���.E(����� :AY�"D1��)^��0_=��|
(�o���(�������v�t�S�/��U
x��v2��S�{RϹ߂XfP!I�S�j�V_�L�?�\YК������!���'���w3z�G��/��H�Tɇ� H�:���>>�	�^�m���BZ,�����2%�~��b��x�P�t&X8З�e�����#6��br�����F���Tj[pܒhZ��|o�{�
��oh_���B�Z�`#�w~�OiP�m����F�[���մd>^��s@$�U�'����k*�ڽ�<��p���G��d���t�7/�����7@��≲T�+\��kj|"�9��Y�G���7�{������i'�E�#��T��瓳����:�^��~1����+�}f5�rC��lq����Z�3 <����������V����5�Z�ߌ�;K�|b��ʒ�N���+�NR ����;Rr���ы�ĚIu�ZI�(���J	����
��qpݳ�3-�`���Ӗqo�}]��`�t���z�������/��_Q��;�{���H�*�UY��y��:�X ���Ba��V��nȷ� �Y�|I'}/E�݀̀Q�;*�/�M�"54:b}-�Z �8M�
%;�D�L��!�������,�5��~���]'�:��?��x٢��J5^^dR���+�i>�����W)$�N�g�r|�	��<�fI�?)S�Q��>nCZ�^1qĕ
��d~-�D�w��\���j���EI%6�E�!��f}����K��:4��.&9,ӕ?���N��'//ǔ�&�Ȥ�0�b̏P��}�8�߹鋜��Fek�f&���W���v���u<�X�x&C(��a�#ڜ&�t�\�;�Xl����{+$N3��MmL/��M�^,N�����6��&~Ȍ+�P�!��D���e�L�f5�`������3a��ԟT=H�%����L�����P1�Ċ��ao#�ӄl`��WZL�c$�+dj�q��=��S���C�����W��2FZWv=H�3ꐝ��[�6����b̌��2\'�ɥ�SO���{��z%V�&SU�_���`ҡ�+ן��I�U�5�t�2{�3�vL�˯�2C-�@�c��\�11�ag&m8�X��q;���ۇŨ��K��~�v(���u_�!�њ��h�F��l� @�w 4f��@��\�����߹��ηՠ�Tӱ�̈A��\�q�I��{��B����=���|�<�a�.�թ�a�#u��DLC���W���u�,p�v��Z$Z?���Ch/��� ��Teˇ"����� _�����/c�$HqȂ^����k/�KT�N��?�Z� �0��7���%i� �^��'Im�z��~1�벇O�w����}Nǰ�%�s$����L9�{�.w��r�[���_+���0����č�	��y����� ��S�
F�(ݯ&k`z^xL��_g�Y)P.OƵC��<�@8�X�`FhD�{�D+�cp*u�GaLM��%pO�m�5:�}|Z9+JƝ�\�R�,o.M��G+0`(-YQ9��es�����9�Y��*��4x��vs�	�ԙF�#Hk������r\z�󥽯槬�h�x��s��KHLӫ�q`�A����a�%�_�3����\J�����s�1�[d������a4���9C����xD�e�"��Y���A�G�p� nߜ)�)& _ƙR���xMN�.HՈ�Ҙ�H9����OuT�A��^nS�	eڍil���֔s��q�L����9hK���b�D�D����S���9~�#8���܏�,@�a0��9�Sb�ׯrE7�7�T'��|]� �~��-��R�9�⡅��@
�i��1��f��棏����p��]�0�/r�joY���3��v���	-b���s6��2]�^��]T�7n�i��ϝ��za�� ~�4��3��+{@tu:)J�.�V(΀���O��!��"%b��TV��{��LN/���n�3���F{u�2_�d��B��%�U�F�Q?��K�^@Iݻ՞�6a>��做]�:��<UL(�D�xk��y��#���>�o���2�R�2�$�j�dx��hO��4e������
-H<� ����^�6�|��%���8P �{W���K�ᙻ0��U[#C2�IO��3�9�n��b������,���KE����«��;��`�C=\HFՙh]1�9?j��|�:3aC\AO���y����۰�LU@�u$ jG� o�N��5����x�c���-m�W�zqA�6���1���Zy��gf<�D��o~�d�2pV
&=�~�5.�T��`{,�}���n�Cp	��:V�un�7%�<>���%���#�J	��{�=�	��m^��Cޥ&;@:B�1^q&���>���Oy���q��_��B:��˹:�6(u�����js>X!en�j3fȼ��A��uz$�bz"�ej2�P���.H�������d4�a���4uK���-��f�0'�X��Be�+#|����l<��y�+f�����̭�V�	�M�sPȱmU�&T�'ӛ6�4t<*_�BC�]���>���snq�M+����K2����n-bz�8PeFα����e)�`��D+;z���j���ɛ:ؚ#
Ι��ặ�N���W�2��H�V@�J)�c��"r�?����3�>�ȶ�6��L�-�:0$@�-L�*�#�hO���uRq��G�I�6ؓ*.&T�p��I�Ґ���_M��������\�F���h[�G`�=Օ�^�����5n���?!E�uAXdO�5,�3����ԟ�gs�C���T�Jȿ���j3L?K ���4�o��Jd!@�?2?TYN@�HU�bi	ݗ��Q��Fi]�����e�:�>%gTX�T�~D�� <�N�_i�a��n��B/7�waE�i_��l	oMh�xԿ��_g��qX������S1�Md*[��p�=�	��jg]�,�P;���RMs�dqb������a��\��f3M��X���Q@��d'��U�3��(�ݺ��c������/L�G%���ۺ�&0l�V!8UK4��75M�4��V�e���5����Wr������I�L�-y:^�̙p�]�Ƅ~���@,<L%_�0��o�Ԧm��x��SؼزP�+-T��Zb�cO�!	��h�+��9�j���Bil3g={�}K �Ώ��m��]J�&�Vom��K�k��v�|��Z�2���@d�+�tպ�R�,�ߘke#��� �f�+�7���_{K�
�2��-e����E�4%�x���n�1YB�Q�J�i�je�u��f�N��{�饃����?�_���Ƃ��	m_���ѫ�� �f����R�=�&�A�l��3{C�%��)J��4�H[��B; ��W��d$Jc�#�l�Ϣ�'(ҬVm��g��7͆�b֘�#��laOzD��-D-��As��N�Qg���j�EO�������7kθE��t�������Қ-Sv�/��)MM6��7���5��s�40��-��:��"׻�m쓰֎K5g���zM
�Bb�r�щ�����Z0x���ߢ=VK�º�1A�:D��h�ፆTk��6����Ђ�륫Ԁ=ZjF��YcH)� �k*s���X�M�S$��my��䬨���a��_K��Τ�9���9�G��b� tC'F�!�<ֵ��|6�Y[[��N:ν�;��0�2Ƿ�xC�O���E��]����|��EW]{�o��$B?1���Mn�d��&x�ϗ�b��S�`���+��V_ǜr Yf���m��.{�}z(�~K�����ͼ۽/H�6d�m��X�(}�3�? ���E�\ \�a n�E�����m�Ö�!=T��WWZ9�	��¬�6�3b�f�A�$
ܒ���p��}A�&�� �s���"�X��r�+-�To8"Y��M_*��U|�� �5h9 ��^���d�F�7��9��:\.u� _��Z ԁ���n��n��M�ųW�|�.IH2>q�T������
8�oh*p�pK��\\9� �k6A���T�B,��&Ϙ=R�#�^�]��I� �%E���p��+�ne��fd~�%Y��3���-������Y�Sx��p]9�"I{Tه+�?~'sw�(�^M0� 2��|u�%F3�~FL.s�(7��i��S
~��C�/�ĕ�R�N�E�0�jk΀�I�����4`�}&Q�-H�bM�c�5O��z�I�qα��rC�!��ɮ���[P�wi�-��_(��('着1��s���gt�)N�k6$��/�>ط��u�����>�W��p�/+��Q�Ao�!�D�{1a�;�f�5�&�T6��E�yM��p�[��t7j��H�wN.࢕�1���m\ 0tÛ8n����"��;.����;~�ڒ\A��@aH����8X%�"O����Ĳ�*���q�>��;@���2�d�8o�O�
E��Nm:�u��'�?%t�����'!��s�7]֢�t@y"�~��ڤ�9�~k�QW�_�t�m�3��j�����*���%�p�5lO�P��=��H����M�(p�(�NdEs�zb��'t�����?(��5��kF��27�<ԫ0@�dN�.�Œ`�m b0�%6R�d�o����P�ۮ��c�=�,9$���m�ʪ;�^vJu��>�8H�<]� �v�  '�W�g�cN�؁W��2\ĩ���@��Gx{S�ϮWE�u��Ρ_ �]�]��W>�(�I����W���үY�"4R��*��5$�4!,p�j���C�n�\p�-�T��۬�3��"g���LqX8�K�w����h�\n�͖��d��A�~��B>�����u�=�ӽX����s)u�M:ӹ*O�`��&�����d��Χ�����zJ;�5���ϳy�s�P��k�,1�,w3�F�&�A{oTz�7aC@S�����$�cxs!S���x�$_6�Z&���sE�p��<���S��0�l:ڮЋ�l���uT��M�}Q�aW�aTZ�lX���¶�
ׁҟ�9I'�j�oo՟��D�'9]Q�HZ2Π%5�� rdn
��nǁ]��U�F�Z/����}ǫ-�G��웛�;�-/9o�Vs�����-���.F��(-&t�X���@��T��T��y����V�d�ߟ�{�'z	�B��αe��0��z�ر�V�ß��B[b<��A���x��)�p��x3��C�hh�D��k/��^r��У^����L]����^�b���z)�I�A���Y.륹g.�*��֕aD��u0Y�#s|3 v=���0�v�t������l���hb��#%ޅM`�hc͡2�2�	��))�j��5����j�P^P�d$l�=u:��AQ�Ёy(�m�����],�� 7X�����~��4��!�ﰬ�B�;n Fiɖ�8t�1��� ���V���Ā��l�_ptR�_�`r1m�M�b����
<R:�����M<�����I!&.�f�����axɕ�,Af+[<땬��.�d��h�tx��1rOI��#��K�\ɧ�E����z�F�I�
.\�	����c�=܊G�	?&�;/L��_�ǌS�[C0�^=_Z&��h�kf�Xem�n� K�G�W Doi����A��v[W� �ws?5Г0�hZ��̊-аf�G�w��'C4y{mS�8��{�<N�T�d�P���7���Zd�x5(�r�DfB}��b��z���:�+T��Z����R��mA�v1e��C1;&/�R:�����8�
/N��!�ȹK�TT^#��E��<�r�}�z�H*l$ɞ�aw҅��{�*Y�5)A��f���k�~R�}6_�g"՘�"vI�9���g�°+rە���>ҰD\�SrD����H9��@~g�_,��B��-+`�d+����t�C�ɉE��^����)>S��|�&K��dKN����!�f�1�:���`Y�?Rn��Z�K��;�Z3b����������o�Ґ�2�_�hԔ d�܃�k�&� ���f���{������H�6%���R��ܪ�\=���������f92{��h���|g1� e�2c�cH�Vp����	G.�rTR/�N�(_�sc�H64-E7"�I�X�!�N�mƃ�ϓ�H�&���'"�`X[��Y�ؚ�N㌨�bUE���E�[��ri����L������v���B�L�N;3�g�p��ڭ�:���!g]{�j6���jM4l�u�d�q�oS\���8Q�m��W
���O괛��n�����?�p��T�Ty̭f�e���&��A�*�B���C�-`!� �&Nd4��6/��=�������W��_�ޔ�4�xo�l��&�,{3� -Z�?��Y8��4b\��1UŞE)}K}�����# w�������aB��L�������$�y`E��*���	/6�A�!Q�����%`�M٧�9��yZ�X������k�k(c;�	W�G|�%�1���sBv���a��N�SM��&��{���r-r$�dRN! �tuE��SO�0ms>䢡1#a�r�
>�
�!H��4��Yˡ,nGA�C�`�����A 	_A�HϬ5�`��p�H]ȧ�x���ǵ +��ʠ���.;-e���=e�,�	ё�"n�OQ�>�{���JtE0�KCҐ�5!��O@q��s����0Rߠ_Sa�	<͈������PmZ�H���%8}r�Sl��H�l�K��W����:F 5��(c��_� �.�ޝ�ML���~��Z�Y�t�]���,�xH���|�3Ɋ�o�ֺe@#تV��#.��T�U�G��L)a����.�Hf�0w|"�9��<I4�9'�?8R�� p�a�/.�)�xM�M�gg��2�riNR@��R|ݳ�J�Y7�ux��e����u���+�7�l�U_��J���V�U�~����N��H�GP�$�926�̈���8��x(����b��WU�����0����F�[�<��X�]T������[�a��r�jE�e����W���(V�}?8$��>��H�:_\��v4aM�Fϭ�B����w�"���Lҫ�,+�ֺy�5���F�0Ɯ)�p�13@��^S�\��T{;�	]��,�;g}Et���Gi�g�O�.���!Lt��_�Y�NƝ���b�q�o�rQ�0���H�E��~�_{�~=1h�T���іma�f��`�BďF�f�CkE������Rװ��S�Ya�a	$���g���4�W!�wT�] 	��X�(���3��i�1R83������T�50�k�����\%/J����KB���O��6��t6��_��G_��J�e��+�0ź���r��wbBrF����A�%�m��k��D�E����$��ىe{;�!}B��̵u'��+�f�,|�e�8�.�U��cĉ���m�-���᷷�-@�����[��?�/�0c=�P�P���#q�e��+@r�59�5h�
���F��/��y��~,zMS��l��-��z=�0'������\��=C��o����U7�p`jR���ܜ� �1�����&&����������<#��`\��3�����w�zۼ"����d��&���ԼrW�A�j9r"�V�f@�x��|[$,��݃7�AN�u�����6� ¹�{�~�!��2���	��.��w^1Z% �Kֳ��1�I/C���?_B3�(����S�e��k(���>dF��"2�^Fwr-	�e.�l 8�6%�/*%rV���y~��0]0���萨�z�Y�NA��.�T����L:�{4�Z�&n?3ە�4p��-�$E8��ԟH�6�!����뀒�>���9@)�w�����8�G��w�T��PD��A����%�6xJĽ�2 �y@�$���O��P,ԋ���.��.��������ˮ*�,�p	
��R-���a�ue��{>s+�ZaRD��V���3��p���fn����Rg����r�mc&d�u�x��j����G@�ۮ�A^g���KF���x��)�+7�N��E�8�3M��LX\�`���F�
�=.�gj#F���(�$
Axm���}�D����w����eJ@�6� ��ԙZ��u.��A�|&�L}����X��Krv�*����]e�\�ɂ�>j���^��.�����T�J�f��#-���^I�O�oƏ�	�����Q�r-c$1��y�1���"��\�t��:�cXh*�o�i�u��䕍�����I�;��5�a����f$ڝ��t��I��t��h����.쒧V�Y�;kS\�4?�c��O�׭��2�xS�>W�('�Z+�==Q"���:�j7�3�.��^���A3
��<���0��؉I V8�D�e#���Q��~��mWTf��Ⱥ�A�2������0��!wf�Ӛ~>R��VB��[,3:�3s&����D���,����:Y��e���g������	tw���C�^771���ꢴ�P��>q~~.ij�w�Jͮ���vһ�I_L�qƒcZT��"F�gr�о��gF�F�O!���� {��ղk�gP"�N�������2n���$��5���ݓ�u��'s�~�����g���m��to��,��,�Wm(��n�S��v����a���,�*���p�jDkT\j2��Xϳ"D�q���􍀈�������� �H�
�2�C��W��j��t���=x�!�e:�Zr���H^חѣCJ�˶���~����h��"G���ϕ���`w:�Zif�EwN�2�;�[��6�y$3�<Co>�b��3'�E"$T}}���ac���θ̪�k)������A����{���R���~�����@�C�_��m�r�8�!�WC�:��{3`��XT����M�\���"���eۯ��*�H�Q#k��o��a{�{��Q|�J�P�Z�x�s��o�e�i��4R�D���r%�rƃ:�^ڴZ�{P��E�L�J�3�w����u����b�m��bp�� 3&��p��~T�[<���?��`:�NM0aT{�.B�-��|'�u��la_h�Y�P�MO.�^������뉷��uW(�Kc�f�lе4:b�;�l�5	�[�]% ���7N�RI)�����l�		����*&�s�Ġ�h����TJ�_�K>�̞p��P]&��0�r��u���Ƥ)7�7Ƙ(����K��6�<�ۑ�t�bm�QQf���O�$�q�s�¡t�_��(��%���w��!�xG⒛��q9Űs�&��̀ދn���|�8.cծ��)���I��G<��w]\E�- f����\�ͽ�c���C�!����6�GW�G��&�L�A �wq���Y�"zى�6�r��y��
߆�c�&+�\�C�W�8W~�rp��&��I��EG�7~?��.���+&��u�˞=���q�6��$Ӭiü'a�V�^��pl?�jz ���jt�S���/V�
q��(��N���=���Z��\aWgV��Л��8��4���%��DC�����,!Z��$~zB�ҽ�თ,f�,`���x���9�l5|�S����(��CKQea9��	:�_�H1��ZeY���NM;뒋�Q��Qf�+Esd��17��ۏ��Wȹ1_�W��%�a��y�/}�%����B��I�FX��6�'��o��,��V�{����:$�0-� �.KA��>�C����xc��V����Fp/�0V�m t�W�E�?b)�8y8�~R��(���'�|��
�q#�;��/J�G3����k��1d17%v��{{S���B��B��"�k��BO~�5��T�����J��MQ��T�I�>6�����+���&���)�ϒW)Uy�6�[$�(��÷%g˵�s
�^A����s�Ur�q��JA�jX�/�w���*[:�t�n���X,������"Q�4���sa�b�Q��b��X�LɌ����.Ƹ��Cw�)��?^���Jo��˳ۿK��>��&��[_�nY��I>�]H�鬲~�������v��M��y�u���^x�JP���+�7��a��۶F�^��
ᦸ��N]j��d�D�☐R����͵d)7<�l�2f#0:I��J�Xco��d�.�X�PY�p!�}�.��a����>Q���k�kͿ�� a��eT<�
	�]7<�B?A��A^ڔ(&t���s�߯]*�zV��[UR�a_Օ��`l�X)�����To!+&$Lŀ��CIUΩ�0���	��B�FGq�-�_m�=��̔�����[:������xԍw�)V�ު�z������I�hR?iX���c|�/�XYp�z����g�rF�mJ���Do]�:{��cB�U潗�.MQ��e���X.nw���$����w��z�r�1��Z/�Y�h�ȋ��{ue�B<*��Y�eI9��&7���O�O�3C�w}��J9�t_"��
\w� �4�uE�/@�M���k���M����wL�3�3��J͗)Y�Q�]�&�c&htL�A7^d���j�X��gJ��p�����B���l�M7V�>	3���O*9}?*��ɣf�謠��K��M[�����_^�ܙt3�*�R��Ք�6T�Ĉ��p���+�w�ơ��Dk�ˣZ��@0��[�+L��O�fK%$?��;�,#n⽼_{eL�wm)x����R�f�[�� R-K��4I��U�da��0���Y���[ܬ���8T��-��U�.�^����2X����\m�l�OdI����x)����V��v�{)y��\=mg���I�<Ôg�|���MD�C��$�XY�B>i~�Y�Eh��o��98��I�b<�����<�dJ�t���Y�5�Ņo2��OS{��$v<�0�5;Z����5=b��6�W�i2��pfD�a�P���N��jdl�%� U���m��v���.�+j�_V[թ�@#���>��	���mp2����V��%~��L"�%E��ulaU��j�w�72��Vy�k�,V����=�H����/���N!񨂔�܎�z�+����
�~�@q:H��ۓ$�T�6A)����ɭ1�"�M�_M�>�-��\��\��~��#�t%R��#��	氌�ӕ�UE>��I��?��7�Y�oލUC��O�@�.��2����#�]�z�T�m�!;c=�i*2���@��8�̓�� ��dq1��A	k�s�H�â���Q䙒Ovra�0�y�&c��C;�O3��@���-U��o����ݤ�"���O�CQ���
�L�y�kH<<��'>ՑS���d�{"���q�+홧P4��d��p)×��1��ъ'|��� �kjU����)� ��;��R\��Hz#����e�EqTy���q���8n�A5�	��,�/���T�3�V89��=���P�f*.��$��('.�Ǟ�]��9`��z�_bk�{�vcn�`]�}D#I�h�I�GiY�P��u�����8g8G<5�Y��7�+���B:�P�M�x�g8�~ћY�}H����o�%[��r.�ݵt��|h��$n1Nk�8+���%�^?��8���c��<��V�b��[��O%�`�F��@3fA'��a��=9ً��^��*�IΖU(4s��a;}0>�C���r�1bn����Y�xA��{,��*�rn��M��J�rJ�^o&ݰ
�xs���Z��8�ӿ���궀%3_0�Va�hb'|)�����hb�@]���Ό�{]�,�+F�E)Ҹ�D��n��9�8�]�CI�uK$��!�ˮ�>�܊�L����(�V4yV(u1u{��ۉ�x�����i!���3�$.[ڱ�_,��w`BE9��s�����߶�)*���� �4{���?+!����F1Q[��[�)��r�E�\�U�7���k�"�(��T~�ݹҏ��t��
4ݮ����#atc���^�ݭ������m<*�����b��Y��_��W,�|K���&o m���ByO��{�H+g��pg�5�Z3V{Nc�5<��9��"��?���{%W�p�F8�o����a>	u�:����]��g�	R�<茲�txa�j�!�S���߅z�]b{��Ӥ��??�3~���N�٫15���ê'o��q2��K&q��]�{Z���(/��~9�4R>�d��^wѵ�<�E�#@̼}>e���J4�ɗ$O���X�Al��7�F��W[�������Z��٦���,����էj�q[3B��7 h��-�b��l9vx�)QLB�XsQWH��B1In��3ͥ�!��hBI���y��d���]�Md4z���١�n�����3��i6_��z�!ˏ�^��[�>�&'k,��t�c���>[���5�,����V�������a�j)��� 74YA8��D�D
�{�h�څ�`��z|P�GX.�'G*�����X�C�'���-a��T|b/��dz�侫�J��p�t��Pg�����4�!sSy%�N�	}�]�_\
v�ڷuI��K�3�܃�J�QY~Q5��ff"�=G����;!���`Y�H���JxJ��^ÕމIf�g�ũ����o��4��g��P=Y-/㉬|�^+,~yH�}X_Pu3rV��0h)�W�e���i6'7Z\cڇ�c���xcش��(�ԭ	�L.�ZWb]���X�=�s�b�"�7 MJ��>���6�d�h�"��NG7�0N��X��6��r"Wx�Y�N���T@x��}� N�]���vJa�44�����q�{��>7��$��R	q�� -E����|��b$�_(�st 'N�l�2�1�#4܎�u�;�]Z'2b���R����2]|&��=��A���h�|�Z�����(�Qo��>����/8y����Z_�~)e�:Lj��v�oْ{�Gݙ��8�̄��
�v��
 ����V|�#���-��f�1
�g�
�\��;xPݽ��P��@�����ʋ�-���VM�|2-hSI�]��|!�fl�i
<���ӳr�N�m�� bm���X��Ã�rM�Q^�f=��b��nI���HLOJz�U��It<�G�ֺ��QH������z�����53r�]��U�/'�'��M�k�aC�|��A�j�G�kLѰw>aV3�01���K�tSL+|�zW�[(�+h1���p~tJO�+���m�JH�h($g5�\}�Ϊ}��RɱN�׿���B4[]몈n��T����V|�?����3`J���[����p�%IQ�F����T����H}�.V���}r x���RW��2����.��K��u$����T� ��|�	��*�߸F�X��^ԧLo9����K{"*�������2�B�Y����,:��(�n �&��-�:�z3"�jR���E�>=o�$�b9%x(ԉ�M	���ẹ�G-�`���ߓ��P0�K*�\v}�|p����,���ɞ��kYѮ��< �o�il *Ks"Q��"U��_`�IP8�FR:@�:�S������aqK"Ƴ�(jT����Mu����u�i��<�=�Y1�u�iW��f�ra+���}�-_F?K���kJpؾs f�Q���$Jp��%BJ�խ���4���-:v��P������F��Q����~�U�� ���0�~�z�D�8n�~�����d�c/n��;�c@:���'C��.�z'�O�y�	�����̫+(�o��'��Q����q�C�QA���Z�ev{UQ50@:Q��/_���}�i�&��wN�-�A�kM�w��y�CĦ�-P{����σW�4R ���|�]�����O�]V��3!�Un�'�9�<lAR�Q�{g����s��c�s�Y��>	�W��쑱'H+N��O�}�X���W�4UY��O7��n.��]�ƫ������0���P4��60�������߄c;�[�Pq�%m��x�	��!p���y?^k��iW�t������%lE1�僯L���D���#�&�]3&�1��A�1�����IZ��?0Yc!�H��b� ���mNw�������/^�+�K�G��[�jV��LG5��ղsk�3���O
h�)�<Z�D�ZyA��ʀ���`���HJ������2�7�Y���[}Ō���s�A!�e޼��$p$·a�D�.���~U8j�Ɏ��`
ubP�����*Qc�C,�D���5%�������K��żt}�I�����s�S�����7����:�i*�\���	�-B��<�L�5b���$�h/�c��/wR�C�t(���je��!���;3 �`�M6MeU`T�`�@�V�zV��
��	�T���"��=#�%	������s���W
}�v?�,������cG�?e�&�9�ɔ����v5^�*声b�|)x��t�gU'/��5s6-na9�jd@�s^��F�P�B�ф��u���A4��GK��'��'����Ӻ��gC�=s��A}^�h�:${���#�����%�+RU�G��5���A��8�����W7���;J|÷媧���n9�v����Va�:tEW�3e�IR.�;f�q���:�U�T*���,r�k%8���{�w��@����F
\`"�m�_pf�c.� [�+��s4¹�ۨ:A�U����o�!�&�K�~|{)H�x���L9yT�	�p�����'Ǳ��K"�9Ɓ�
G܌����-��?��~^��~�J�H�z+*ԃJ�N���Nj�-K����E͇���q�a3ɽ%ub(Ȟ_Qo\��.�q�sś`�D��c����b��
<�E��[+���[^L.��F%� A��}F���9owX"5<����k�
|H���*��u�JW���V�k���������g9Ȼ e���?�&�_ϐ�<� \W3Dy�g4���l
hD�Q��e{��g��*�1&�(|����n%"�9�K�џU���|E���g֪U�Ĺ�[��Ʋ�R��Q����D�v���F�N�2�~��;g�K��f���ri�Dg��1�ڴh���K�H��LӨѰ_8tD�������Jw?�­Q����M��u���o{��~�v5�������6w���ԦQ�l�z�Bo(JRaz�`g5�|Т�S��U�C����Њ��!��뚖%@D��I��L1����~P�l	�šx�c�e��ƣ�r����H�Ä�5�c� ��;�O1��yQ+�Y�Efь�S\��}xŝ��&��r�O�B�xL�d�{��|q��'T}v�5� �K�>B�ٜ��׉b��g�MSO@p���Jm4!?��,&���<��P��V�h�
���<NY[)з�O��8�7�����GǝI&�3gN��d9�ӿq�`*j�s���E�/�=��nR`'I>N=6J��K������U>�R���(�E�$s����ɡȍmYe� �ϴ��q�d�e�@B�y�J,�ns��g�����ڑV��p�LZ&>�гb���ue�_��$-�o�gcͨ���{�Q�}��,\TX<�=E��&�vН����5>�/@�㦳N�)<N�i{��;����{tP�ɾtזpc��|o&����SA*��������
����'釒�5�
�z��l��ĐZZ�����B��o%����Hs���������� �gjކ��f��
���##,������4g�X� Z�q��{F�������.�'Y-6[��X1�
Ҏ9����Ӯjz�OE^!�m�f(X��J�\�m~�e8�I�S��I�J>�?��qJ�B�z~�T����J�8�9v��[�N5a��|��@k�v�/��$ޠ[Puj}V�iB�Z�eb��r��=��z�o��(CmOßrH���wZnE�8��J������\'W�ˤ��"l��e	Аם#�nͤ"j�\)-���\Xu�(؁Q��#���~8#��.��eQ�\�d��G��fx>��Z{yq���':	D��/ �#N�ɧ���9���w�e�j�2\P)W����'�����PuO�=��!s����`��/�s�!.��He��^uJnyw�X�\�Pgm4�"P)b\�^�\GA �28#��4q?�T-+<�i��4+�\{�~�]�+y Þu��<�L�^k��o��,
/�~�Ss����̺e3[#'=p�aަ�˻����*�OU(��� p�?�T����S�J�Y�w�8��5��eU��uP�ϊ_Yw~���$���$n��Ig��^��J#.�H�.��a����������`�[�}ǔ�5�x|Y�J�Ώp�H�o� O�ij��⑮����c�iŮW��m������Ͻ��	'r;Y�%��uf�T�T��Y�A��n�����]�w����ܘ�Ce#�v��d��>�J��2�	��g֕���Զ�.�"gqq	v�/l }��"P�.w4`e+���U<<�]U�N�����k$}�%��қ��T�G�1,odV�t���Q����=���nӎiI7��R�zb^�s���*7���s��X/�;�R���~�t��?�!���������qZ+b��$��|���`�k��b$�	3�6`48��֑s��V��`nZ�l��~ �fy��>\1�+����ȳ�Ҡ�TV�1��1s��	�ޛ�&ΐ�<�A:�"�����;��
�ᄋ{5�R���^���-�=�rF�B/s�p����"_�5`�;غ�u< �zVΒv��\���э�,k*ɷ�ϊ�x�B��؎}�$�&-=#���J������p�R��%R]�z"����l�]�x:M#��7��	��wU��,��OF	˖�E�,7��,��ms�դy����៼�@^.�C���p�6�;�,<�1���'��d%�\9�Fҿ���4es�j��-w�!�c�ьR��O�d!�>L��s��ʖ�Yð��t�� c���k�|S�F?��BP`����˭f����~�	��Zw'��<%-����2É~h2IF�衜�HڄD�$�gP'L���=���!Y��Yt�G�9Z"p6�#����
]{�����϶|;l�Ga��
�̣�����٬��Q��2�����pITD|F0¶ s]۝�a�o�BD@{���u?���j���~�i�A/_A���k�J)��/B�E)<�~�!�k��pg�B���Gd��"mS�k	z�=���t��� T��j��Q�p[��e��9�L�^��}��4{��,^�?Ρj/Cnq�� �8s~�N�C0}�)R�5�H�����韶�>�2w'��v���>u��
|m��s@VWh?��Aro��='Ry�#�Ep�H���<>wW�D&��!�˰/���� �c�]�c��`�9k��ź�=�֫��v~뜜�����b����a��:S3��#���_Fۢ(L�rA+Wm'�_-�/�)l<J�{A������Nl�p�S�"�T�RK%��]ձLG�j~з[�� �vR	�KAo� m���v(AS���eC�����T�i5Q|�Sv1�M��;P�9��Z�rJ$�'�y����� �`�<�"Qb�	:�g�>NP8���I�}KCW�lmڃ3-J�h��%�0���VP	f�=C���zi�5��������������ƿ�_|9���t�.�,	U���`h4 �˸��{O7�\�E �����t�x�1L���U�,O���~�lh�TB��(��N��u.�@���G]�Rh�旃BC�
i�V1�X����%Sx�yQm^�"�*`,��m�;1��5%9��%á��֧�|'�b�*��] g<�j[�.vV�H��*G3A��#�g�ћ�&#tV<�s�.�	q� Yf;�Ì�zCZea���{���]%�fY��T����1����067�"#s�# ��j��K̜���]�C̵m��.�L���IX���e`�<�&Iy}�E�a�aE�ݻ����@4�d�EI�' �F8o3��I��o=Ĥ�;�/��&�2V'J�Z!�I��f��|%��_�8��1�g0O�C�+��[��K���p�CK,-T��a��<����9�I��F�J�k�ȿR�D��I���m�opr�������
���CD=ջd���N����&�s?޿�5%��X�����p������d�:�bĝ�$�s��Y-��ϥΛ�HH&��LȽ�&cD߀^��O��hK_E6PZ�uk �B|?;G�O��|
��ֳ<�C��s��KaLgE��'(�2//,)�Ⱥ��<� cw�a�u=w�p�[�8>=E�K� C�I����<���{Mr�4ԯOa�|��**Oru���?D��ɔ�����M���fa��,g��'���ܲ�&�F$[:rI��}A��g䉄x)�w,$f�X�3N/�n׹ߒ�"�{,_؁qo�r)����c������
-�Շ6՚� �wS��b��]67m:����{��|St�F_h�u;_v��}��9I���{sb�P�����o�$`d8
:�F�H`��#U
����`)ߦ^o����5�����^8���9�޼�7�h��V���<~+��|���;���}��2�<[ZZ|4؋�+Ӄ0�oaqk�@�a�+�H";�=l��!��������`9�j[��/��l����3�;&�������g���$� 3枪y�jt�����<b�Z�0��m��F�1T��+���e��v3��^,����h�\ҟ�4}E�eA7�M�Ʋez�q�f0E�d��/�s�E��S��EN�# LU8Z�����`K��%N��!rpí�˫���;�C~ɷc-��EC��0��8����_�� $�"�D��I�5H'u�R.ȗ�7�h��c�"��f�/64�}Jit9:��,Wv|�I�d@&ƚ��q�� �yC�EOND�'&�)��O(��"��	s)+7Wu�p.�N�T7=��H��ʲ��d��ܟY�|zz�vQ�[ȴ ެ�b�Wq�a���ӓ~@��D���l+	�d��S�o���)3��z�C�ҟfi�]]���f��b�߼��{�&TnN���q��z�h#��Q�����39�J�� KWd�+�$X��ISkbmr�)�(2�%��7�ױm�0|���NjB��� ��+���ú��̂,e���]����L�Xӹk]����,q�?������������hF��R窩��{�#:�U��߲�<�����z?�I!�**&;5K��欖���^�y��b��	���	:�vC���}�&���[:�\V�5�V���	������}o;+#��&��_ց����t�H7�}��}�;I@�2��[M)3~!��'�4�X�����&|n�Hʫ�T2�sI�)U�c��k�s������y��2|%^8�#bz�r�h�@��0�U�>7 ?CU�e��}P�t>YR�n�~�kl�g�.+r�?wR�%�?J9��(a���q�m����g�9S�� �K�㴁����}Q�P��?������Q���l�꼙gp�T��!�������A8��a��0۞#�f�,��Y����}�k�+J�f��ձ���W�7�҈B]���x&�� Gx���uKx���&9m$�����8t�N"�l�I�K'A�Q�]P��(@����~�"��!���U�Y�ݹ�.��J}�s���k���w�%s�S�ڡ��g�{����X������o�����Q�\��5D4�|���Ϲ􎀞T�(~ ���|?�kTIٮ�+E��fH�O�Z�E��x�m;��Zjک�9iM'�H���F�}�hMtw	��n��\��Q8�����u����k}��G:��C2�[�GV��]����l�s]=5i�\�i�rK�/��P'�gT�Ե��0z��v�z��?�J�d�Է�q��Q��?]+u�O&�/!���T���X�P��F��8����R��gh�(#��=<$����ƾ0z��>/�J�*����F�]}��#�hz����~rb�����ᚄ�	�wҕ�|���GA&Zce�|�W�eLfXǥ3��yQ��x�S�����-	n�����_�5���\�����z/�@6�KcL�*�@vQ�x�8���-$��")�b��VM���]��V�	�6�V�%���,�`��t߶�e�]e���2-	���F�R�
,A 0`.�p�%D��1���R)70����+r���w[��[^�d���s=� /�j=B�5�s�T.=+B�6_��3��^F?J��)`���ݚ��Y��JC���/5� o-�Pep�=[T% �;a�]f�K�U#R�uB�,)7 ����}yc�8����{eX=��Y(y J`�g��xQ��q�:nkݦ��$c����*B�m���]l9��`��y|�I/�硿���(a���giۼ���
�|��P������>�C(/���9:�����.�Q���-/��τ�<���b�)b	qr,�D1�>W,�X3k��e��}/fn�h���J���*;������	�+�����U��]����S��8k�Ѳs��WW0hs���Z�.ȸ�ʏ�%�g��3P~H������S��Lu!�T�kF��m�P����,oߙݦ2�{c�a���s����0Ա\�(m}M%Z�|+��9�ؚboȃ�ن��=�?L�Uy7�B�cdm��cd^U�5
4���f���3�.��0�/*Y$��u�iWT@�>�j=`N�w���
D��a%j���
�#�)�[���zĠA��eI����V3w� ���-�1Hq�Zvf��x���Us<���������A]om�.:���ՔQ����J���l�jof�x� �S�3�	=xy�K p�tǃ_�Aح�F}���+ܻj3�������i,��dԄIP�ޭ�1�5��? �П��7�F=#�8f���]�Qj�~/G+;��NU�Z]x�'�˦�jxȴa=�Q� ��2J��~�z��%L%v�!Z����E^+�K{�ûKWC^JR�HF��
Xxm�ɜ`��~#0"L���mJ�%����)�]v�!lB��<`}f�p������C����C�2�ɿ>�ߎ�>~�X�5�J�K&� ����/u���Ej|b�__,Պ�j��(��1m{��]��KzXɌֹ	 EŹ-d��':���MՊ���������`�.#�D%��5�𱴧v�W�4C"]G�O��Ǒ�����3�� Lx�yͶ��8t�u# sj����|ǭ���++�2^�o��r�	����{Rq��H*"f^Y\��=�˞V���u��;ﳃ��~La��E6;���}.D+1wPȎ㩯�h�	��:x��;��>~е#�ٖ	ot:v� �3q��׀vR۽�s�u?"6�}�D$��ҕ��@h$]vB�{y��B���Ai� gh}]��`�>�U�S�H,p�U���V�S.\������i��ׄbS�#vi��F�c\J��X��$�$��ˋ�r�����d���0�M��`J�ܲ�u%|���`;�!}K�r�I� ǋ��GݍӔe���U��,�Q��<\�G��Ae�q����.i5�K\��{q�gt(T�s�x���@)BUH�����Ldg.��*�#l�C�aː"�4��iձ��l�]o��)0-sV�"\��6.�pi�#?�w�꾯E��lJ�#��Ǹ�'�,G!@@m���V�wuif����a6D�%~�S3~�dJ��"�kQ���0MvA�We�%S�Ψh�a�F���3~:����~���=�`�&~�{�1����r�/�D����t��kTO�qo��>xk��E��A�Ah}Pmg�=v�Z�e�i<��� 1���2H*=�KA�w�o�j9Kɲ�b�Ϸ���u��7���ۗ���1�C��pIe^Z��^���\��}�)�M���n�FEF`P��l���30g1�M�
�ھE��ۭFOȧ��j~�ݒ�ytG����c[߮r�ݒD�V����&[�;V]��w$P��m="�M׏ѐ4�4A��Ұ��U��*]9(';2�i~�v�Z�hH4.�Jfk��`-�N�����t\�u�aaPV[��ۛ�)̠��<��	���肘ڶ�W�Zu8�"� �|p_�&.S�В�\����|�� 2�Qw��G��֒�UD䒷ʹ��� ��_����3����Y��/Ƙ��/���8����g�ܗ��!/)��U�Q��9s��Nh�|(�8�΃q������'���m��4S;�"�c��#��/zf��>v-�cb�1@�+�j��4#'�)qI!�h��������*31N+rN�g�ǭ[��T'����\���!ь��M�-2�I�	��r��3#�$G�M�TO$E�tכKP����#CG��~����J�ް���g�S
�����FgH=��@�ɺ��V�v�g��*Ë��Xڷ�'Y�+����3��}
Ms�ܶ�l��(�Ƥ@��2K�d��[��w	G��턓��8�ۣ�!�qcd:B֯t����c/�mq�g��Ho+G�"��8��ݯ��E�6p��J�)�am�;4 뛢qI��\���h8�!%ߦ����;����˵2X�!�=1�P��Z�bt_��%2�����\��P��Q9׹�$�1ek0i��ӕ�ĥ1f�Sv�$�����!<����̖1�uJɾ{iE���A��c�Q��0��tC�{�G�i�YrJ�)���K��0B�@�Yִ�����~w�CJ��'>�g�ȴ���*+��$�e��n�f= TL�T����>4.	R)x�IX��%9Y=�"e�xj��E�`����_����6ʲ��ק�V�%���K�ϋ�F��mƧ�Ҹ��}O�Z�%�-G�i=��!��Fe��}��z2~e���!ai豰�Ț��AY����Uy�~�g}_\0I=z�����,��ƚ�Q��n|� HY�٠+:3w8��[T�c�w\�G�䅑�o��� �<n�U��"���峳`�n7+H�;�&�׆��O�=lKoZՅL�*s%m6���.G�'��d�>L?~�H��yW�X�x }�ig� 
��w� (�1�ه-�.hͤo/�1 9'�+[[�g>s�Ep&g訸�v=��j�	��_x�B�r���Ω!��$*��!�����!�c��:4% ��s� ���q�t5>J�b�{@�_t�6�P����ֱv�<� ����}�������䉮2]�-�١�7�	��-%4>E�mgk<5�ā6�Tw},�ak���(�ݼŁF�lЃ�sO�Z�6�7S�Sf����b�������*ޢt_|.'���x^�ɼ1
�>�9J����<.��G��!���&�p��#KL�s� �ɕP�؇�/���ޭS(�#����)���@��ȸ}�T#HL.�@�	c`著i$P��a-S�ѻ�X�D��qb�?�3C�����2��}�S��IgD~�`�∨ȉ>�5���/�鳺Q�[d��g/��L/0�$t�:�j:�����u-ޅ , ��_�]Y6��Y���A(L��*�f�W�H1�L8�]�WW�ܵ���	܆"�fJ�Z?'l3r����J��!U@�J�|� h<qF�KH,p���c����4N����b:?
S_�b�H��%�X��e��NC��+yڬh�?�8��b,�8Mh�Di{h��|�`��ײRJk_��٤��tN�AH�D��6v�čȑl^��P?�����ض�ul�C��t�f�IvSG-"4�ĵ�!'k�~p�0nN��zd�G`�=8Pln�ń�4"B��X�ds�u�C��Kn�����TI��q�ߐ���\�I��/����Xk��b�TI�&�Q<@V���i�R�e��$U�� ���U�P{C,�/���H5U��B�����Q�*�7�}?�����Q����M6�ɱ�O��I�Y�X���;��'i�AKG���r!�!و�E��v_���������ɬ��4��F�Q/���/�7�cIt�	�5��W;�n��M���G+i(E�1�"]O��������%�@R�oG!Afs�$JֈB���+:�B�_�x�a8�g�\D�0����y�ѓ�w�&>�Wʝ�����6e���B��{(
W������}�§I���HmE٬w�	��C�f��7�+g߷ �b����o�v���,���(�|�0�C��ߞ���xUL���'���b�Ms�I����?A�VN���3�R<����)�R�.���!=��xi�����K������v!��	�Z���SR~�9�@�����Q[w�L.�-�4��S�3R��Oo%lwT�&�k�O����I�V���@*@R� qC�kVa<G��M�
i����S�Y�.��-�*�S����F��e�NS�>�:ߓ�w�w�:}���F5M�>+�-65�yQ���u�a�=A��6����G*z,e,N�8� �F�pɼ.�r\���)�����o��H�:��H֪������r��h��}"�և�L�$�N���u7��>�}c6�,m���~�Q)�K�z�AL�.N���!�[����}��,��'q�Ɛ��͑�Y�D�^!a�,�<�B���hG�]L釧b7���Q�
��*zm���O,�+���������O\ �"[�tc�ߙSg���xu�Au(u!K^�q[�<[v�R8�U�!�0={�g�M�F�c�C���0��w��H�^xA#�逩Z 4 ��r�ƒ#&�[��s�Y�*2�dյT���dl���|t)R��B�&����+�P�<ƫ� [�R7A�Qr��7P![��|�e?#����>E��g�"�I�w؍��N��ˬ�=|��o�u}�B�4�ų�Z�< 6�&�����Y��8��8��#�5tP��P�,���fg9���V_%��_﬈�Ssw����Ѧw�Оר?\��oq�C�_`O߄z0��6��)qEiz�[u���b�������݀Q\�����7@�.��{]�0��K�pX�o����pUk*�
�J��6#ǒ���Yd*��/���u�|�<"q,uRn���y?*�����􎪝���qҥ���;�<�5 ��B����"ڡD;�����L�O�{p���5��;�X��-0B���l�U�.Z��s{��<׆��r����H�b-l֢3�a�����,�ޝ)����Io���"`�#��Xu�*��:�N�E��([�"�x��M���T�
�-����� ��j�M�������u���-�+FݣX��aLϪx-խlݺ!���T�P٧�& ��g]�)��,x@�Q�sab��6��ѕ�P���$f=�O�f;ma��<Y�����{�٬7���a��ն=q�𬯐�B�
&\d��6�R��DO�򊅓=)*]m�>�ץN�ٯ���EU{[ӡ(�Τ��x ���}&��8�)�o���W3���OX z�D�rY>��L=�*]�hcHDQ俹G�!�h��(�j�pJ�����ת��8��
�E0Y��Tfn��ڱ��ĵ`Ծ7u��i@4�"_��̒?��=��%�A��#��a��t�sy~n��l�Ԗ�#y��g�'�+`��q�$�;k1�ɹ��%=2n���y�	"�����i�W���L{��"�G$�,�eN�R�tr\�ĩٔ�p��<��O⤥����#@"��V�VkuA7�Z��{��ኮة���0�1%�i�(s��}�B�5h�`:Ǩ�_�6�3���M��uCό"cm�_CE��:�KO( Yy��޷�z�B��ڐI �r�ɶ+(pTf��<�P����w�Y3��,�V}��A�uv.C4D�|�%��\�?�0f���cc�
)&S2��c�ma}an|��pK�f��\RM��۴h���Y>VP��ަ��AX���r�}�w�}�T�b#�x9�[�<W�C�d���-ӳ?�t�~�����2��dɣ՘4�A�s��hpa̕���"�ؠ�Giu�ޔ��A�M�ᩞ3r`XF����ţf[q�A�Yd���z��`�a
��}��o^l���'�A'�8����aCI\D4�r�3Љ�/�ŶA�*�ѥ�:/������,��xї��o�JZ�WY�"hOF&�I����x�}�0�:�+�z�� ~Mݤ����+���'�� �`���@b'�(�Y�H=p�����\�s�:�5��tϖ=��]�ϼ����g,xJ�lE0�"����0J��^ͷ����0�L�5��ux���I�d����IH3|z����+����a����
 a��e��I�-w������^�^)j]�D�͊7�	�Jȱ���6T�9Y�hh��2xch��Ֆ����{Z�c�+'ILm3 Pm��_�������!��%�*>ha����e)6� ���8�=cxǊE�W��^da�,��5���E{�)���$�u���㬎r�
f�啫�&jXd v��E����~�ob�6��'�6U�x'�m(u�uO����t���6�>��W��FtR˹�[� D���ƵH��b�hz�R�};@�-�<�\�WV�˱����7P�]��$��MD�]��!��ÞGr�v�@�t ���2�K�8�������9R�<���g�a�迊��Ԝ]��/��o�q���<L�딾�!	����C��'�!4�|�����������z��b-��/��0�8�e�^�D�l;���I�$�R�?֧��CvZ�yd���<��+akr��,u�d�W�{ ЄN4vȀ.7�[�V1�]'h��6:_��:M	Qz�=��g�� 7;\فl��O�|uT����`�{ f���f����ܱJ�_�O70'ZBSq[�ߜ��z}�����ܴ
f7����dH��I`�U�
*��3C.�n��%�C̲�ΰ���D��Do�q޵Dc��7yO|Ĵ��}�,�vz@�G�0\vI��wt�S��%���N�>��~$ϊ�g�3�Ԝ���Jl�#P&�>���P�"��w)�ǧjZJ����68�`�����y���u�h'���[a4'��/S���E�H�{cf�Q�5�kD��1���?�������8g��P7���Azް$V܀J�*�����3=0Ɨ~�xz �/�=׾`�g\�\_M�>����E�g6��.'�`2��5K�o{^�`+�����q5��㘔d01}�0�?�*�2�"9I	�g|vю{v�]�pM�󥹦�}��=���o��ͦo�IB��,y/��3�F�+���˖�ɱ}E�:�.�E����;�p��yd�_m}��"�c���f3&S��d��/S���v�!�{p�B;S�b>"H������-�����Na�y�����'�TLs��	5�z0z�ͳ��a��f�lA�Ը���rW�n����-���kӶ/��3�Vɺa�=��J��.4l�x��{���G�?G��V�9�'I]@�+�Ǯ��Z�W�%���!�:n��&�oH�T�����(��-~�� V`u����g㕔!��f��)F>��������@�����$��Vc��z��W��((�d��;��(L�����,�Ɇ5#���ep=�P���s R�I�.��.��;��I�ac����k�!;=q�$��t��9��tw���B����������I��D��}_���O�L~2���X�ua��MŎUN�h��)018�5���7�m-T�б�[��O	(IΝ�}�$i��k�aJ�*���%gQ�2��`�Ɇ��T��d�/
ƞ}w��03nv�x�-̳ސ"����De��@��iv{�6%/a�!�!8��^�P�z���T�E�w�v�͗�C�N4��Q����uY�$����2��:���)شX�:�|$Ԡ{��=�9}�4#���&g/ѹ	��1�'D��.�B(��W���gg�֊y$x��
]�x�̓|7��<8�-����)�{���zkhh$Ԙ,O|s�����%)��� ������.����y�uVR�	��_H�� ��mF���'4��!Dh�0��Fps�3��>��Ѥf��앞q)�� ����F�;�������l|a�� ����lC����H6������s��z)���`�8�v3F��@�s��Z�3����J���K�.��&�:AO�!y������#!K����bq���C�~v�=˾�;��zF��dJ�s�~�D�p���MM��SGX���] �Ħ�5����U|��̾j�A��f�-W��"����m��F��tǽڀ�����+P���:߸��랎�+���<``}*�fǡCY!�J��G�y�S�a�� r�I;G��u�cA�ȼ�}l����� J�僨|+e�j���t�(q,�!3|�ct�>S;�~)@�L3K�򥨉%��:-�Ji*uX��+�5�{���Gd)��*�町ݒ�\հ��g2��8F��e��w]op��&�*�D>�$c`y�;��=c?�N(�E�v2&�vc��D�yb�$
�'PG��/t��w����p?��>�E@��UR�ܳpp}�L�hFm��g/��G��o�O�Z�گN�y�\�R�A�K� ��My�Z�il�b4|�M�g��5e[Ke=I�[�ИE&s^�P؀ڈ����t�6�>���kߑ��녞�Q�_�N�1�3����&+�x܈Z�H��i���ÓJq$?��^k�i��>�;\��p���8�ދ|�����z��z�m��=������v'���N;�̳�5�A
��;ߤ��Vla�W���L������6-�4h�g�6y"ˊ`L/�����"�1l|�Eͳታ�Z���j�%j�rd^����J	���-��=[������������w�F�Z&�ê�\�h�����<�y�m9{$uy�.
"�[+��7���.��Ao�l��������ˆ%�O��FN�EF��HWko�hh�Q)�~KC�VM/�d�HZ�y�j��W�ZQ�.����:G"�{����C���6�~ُ����ds'i����E��H���j���7}���t�-�Nf�i�Y����v�jL��.,�sI2������Ɓ�5ڣ2�9�T�C
�1H>�0#cPP?�A�r�T�]�N�ơ�{�����zc���>bv�T�&�O,��BS~�j����FxiⲨ����oGd=?r������7�e�f=C�|-�hħdfp�e��KK<Q=�����Ik8\�� �l�T^�ě�E�:���?ZCo,׾m�"��Y�'���$�k�%.��A�@Yܪ����,�K`#.R>dkɬˣ��n�4Ͷ���yt!���d�Yi�| ���FT�U� bǗ�߀8c��1�ᚾ=��s:�9�=d )������J�����e�P��ց�^F�r�y@�t�-ca�-��~�*��1|��p��&<;�pD��ǠIc-r��z�͎�S�VH��(�Z�W��bPT���[�5r��7H�^�a�|���f0�iH!��t��K�zX���:TI���*���?��TI���eW 6��d��U�Aw{��i�"������\��Ш�O	�2ZdE�7�!&:e*|�;6C���@;
@�:���~��	�5�U������Խ�J��90(-�=?����<���?׮��l�+���nɚ�{�S+&X,��X�;6�g_�[�Z4�L�?��Ts�����aS�����?�6�����w3L���~�"s�-k��C��_Jp{>��+�FO��Fl]��|	���dk�ͻZ��%���"M*��Β2��ˤ
dL8d�Y�!~��T�>=y��v��;����_M��ak�Y�@V��BXT��[�bҔ��լ)�lƬ����̸����P)hj�|x"��-���ֽ%����'a�͑3��)	�\<�ڞ���j�;�[>�C����!A�Ґ��R]�"?�V\F��̝������%��V�T�Oz��ޯlz�h��`�vu���p\G�=Ӫ�Q���4
v�[�5�i��5ŏqG\��v��o��h)ޑ�su����O�-b�_��ŵ���Bʹ!*D�%�
w���Zx���H;lb�Wn�&�cl~���$h�
Z�H$"�� �)�D��%PB�!=A˰�����q?\��.?�H��.'���5 R�XM��������Yz�@!W�}�z��F���I{3plZ��t#bT0�U\�x�>1Um�y�J����Y�ԤВ�dv}���m�C\QЖ|�͈�	�o�	p)X�|Q�OG�I�@�MM�y�-��u��L�a�H�|G���`rO-�����vg0y�|��1Q�2� [�NC���?c�N;-�|j�E]�@'�{j�>��k�ڶ|�H�>@ ;�����7HHW�w��U�{t�C*��=��:�9t���!'W.�q�þ8�Mè7Wmhv�$u��X4R� Z9U�Hz�ؿw6�؄W�gG�Ğ�;�T���E�BX�OU����yR��r�̯��3�	�8r��v���x��y�ʹD��;Xli�t��4%�v�Oÿ��)�e�;W)�C^���4���݀��RK�X�N!6�Ϋ(36S�F_U�:H����T@o:B��uЛ>�ݧx���z��H����v�.!��~������"�Q�w��ys�kA��g�anO00�Չ�Q��O���o��T��c���~��5�FI��E�Ǟ��-�a��o[
�����!���n�!܁��Lv].�O?��O<���4x�Q*,w�����_kq�Ddha�^Sp	q-��y�Rt8��w�3��O�m�Tll�-��Ml���mTP��������9�Չ��ݻ����G��c��W�*���Y�{Bd���	��*��D�T��!C���o��ʽo�������G���C�kN��>)Y���� ߺ|}H�p3��u �\����:4O|��Y��Fg�fo�ه�W��y����>t:�5�Tas��4݅�oI��s�T' 2o��j+�P3�e�e�uD���,�-ۉ�X�WzO��{��wFo��U�:9#;�bǃ
�D��ݞ'w9k�u��z~ӥ,���� D�^��w�E�%��[>��uU{���
��@�(��썒�����R���n�Nv=�~W\оA�]�e�Jv��j+2�T���#��T��m��3($"�%�J�-bh댢eb���ݷ�an��������y<Y�`�s�t�۪{�k'�����o���I��#���ZP/K����a���7�]�P)�3��eD�м�g, ��6dN���(��[��l��/qq�	��0vG��7Eh �:��6z ��[f���z�l=�)k5%+�u���|0��Zk`إ���`nj�:�;�6׳�x@$4Y�-;���1Z�h5���m��v�&|?퍡!���ѳ��D����b`ش��{�)��rto�k��A,�2v
��-�r����"����hhhB�MOR7��
ӵ s9^�e`��p���ך~楌>�۷M�#���]����"yt+�(B��n�?6-���;?��^�[�a���S��UV�XV�dQ�rd�����O1�m3]� �KJ���#��<�x"ҲO��EM*��e�h��d�Ʌ D��l�)��d��oC�$e�h.�MuTz��{�����$��WfyM��_	V���M?�H��.��>����z3$-o��̖��Np譵U0+:�ŹE�0e����!;T�#@����O~	���
�f�?�+��A�j�V��������� ��j*�@BCdŖ�;���>N[���@K@�J�{��A�ʥ�=��ހ'��"�������6��XN�Y�іB��IQI�[Ϊ�/C�ۤ>���LQqF��u5i���F�cj�'�>'����q o�����M���C9E�5+�;U��T���Ѵ>���Cf��Z�� ��X�\����=�4}�H�eY�p{�Җ�K*�����G14]2[qVft�B#N��D@�����vX��[*��?&�v���r�NfPO��Ĳ�E�mV熷�q��e�1r�Z�m�a�3�L�������И������(u�鹎%����8tMV�H��W�,/�����Pҽ�$U�d�f*�¸���E����0+ �!��л=:nS,�Q�����{���@�3�-�N�H�"���^v�wa���0w6y#b�qc�(}^���ֿ�u�]��	�k��|Q���Q.6Ml�^�1�~���yC�Fcd��X2(��CK�����t��B��W(���J�^�58v�ms�N?���Y��� Ԥ�����|߯��3����+7n���t���Ó@�*�np�����>�Ig	�����<h�WwF�YPzE^����xWh|���L����Q�S� ^��ӧ�`�h U���"�Чf�g ����
��4.����>��5�$gP����2�2�����_�7�,���֠���e��Cp���T"CZz�|5��������m�r����o7�x��O�ͬ �J��9���
���\1C�O.Zi� �n��&X�˂Q�&�D���ߌg߰�"s��f(����sC_Nڐ{��O��n��R �n�>���ۇ�?$Ni��Ӷ�'0����7� ��d,�>�4�(S�T_v'�������1�-8W1B��i�8+�����]��]m�1��wօ�4H������E�:��,+��D�SL�����O��e�i�����e����x�d3���2��������<
���U����G@p�	t�;��Ѽ�(�UA�s�2i��j��-Ѷ���`��h.���n �)5`��O����<��׫��-�vH�a�қ�/@��6 Ĥ<��e��"�ŵ��w)ϤC�/o����f9&�wJ��0��
*:ǇR8�
͵�;sc�)�A���2A�G)���V�~9�Ϯ�0�ds#0u�c�k�����ߣ*�d�5���
�2��I1�
��5_*�ìR�/+��0X4��¦*Á�4X ��R�{����¼AB��� w�̡��G�r�>�G��k�P�h�+�����ki�EO��R�H�;*��L�>@�׊Z������Є��."]KaMݬ��j�������ּ�=��э�X�k�����܃ŶpZ�$ު�a�ؚ��U�� 	�Wt�3j�~�0�&A�̣ۗ��2�#�V7eR�e5��H2��8A���=*Dv?6s���F�+\��׮GE�b;ǛP��`�4�!U�%ŝ΢ǫC�	2>!;�>W����#ũ����6�ve����lg�.��ަm�
�5&je���=�'�
 �����3г��/%^*E����9L�Va"��X_TH�i��?��{��R��bG�㈴�`�Qh
r� � \�s?�.pF���ґ�3�@�x��� 8����s�9�Df�bō�df�u=�1$	�w07��⎁�2�������aL������>)s�Eyr�,:���h�*|s�t]��4�3`.�L�1MUFx���Ca�X*լ�����o�a�vͤ��M���qM�`!Y�u�dï������-aCa\j!��{�N^i�����7t��bΆ*�RX�8�$���p�5�#T����j,��
%�S�<eh��t�yڹ�;y�w� $T5t��y[*�1x=y�]�UX9^�O�,� _h���}��eo_}C��|K]�C��[��[,�sG؍\G��.�������E&ι���|�3҉@gfz5���z��~�%6��3���@�������*���ȳ��|��Wڱ��WS��}'<|���C�
�"iw� ��H����S�FH��t�(y���W��8��z��/,w�DB޼[(�8�{g����HY&Fि#�p�'�2r<�5��.�E}ڂ�!ph��Q�@ E6�*u?|Vn�1���I��3Ta� S�S��3�[��$�R���Xy$`� �Q=�qGh��Pv��zhSݛ���|bsae�_ jM3> <�E&�?�������ͪG���W$N�ܶL(�lp0�����[���ܩ݇֏�z�ȏ�7Фs62���U���Q+��u��d�ql��W�O�&r�yYaJS5���0�����d�Dɧ��,��P��[�$�ի��k9:��c��鐞F�B���p_]����5@�����>�#�-�[#-5$��Қ�]&-n�M��KA�n�(��=v�9�c"Æ��-a=R!�k�zUšĕ�Uj�����Psz=Ȭ�H5�<��j{��:��f �v+9�NΡ%�"m.��ڍ]���4���S c�4�V��:6(�1��	�.O���G�T������V�pm���Lio(�ģ4���ǖ{T����+�V��Z����SA��ܬ�?ʫ�����k�n(�`�~���T���9p�h�]�Ws��x=�g�
:��!1v?ǔ�g�$+k�\��A�	���#���u�c����#�6�3��<6pTbRd`���۲����f'����s�4�nv�*?[ŖfI��:��ߖ��G-/z�gp5�'��%ț�ʉ��bv���爏c��Ղ-�N��Z��E��}�a�1�#�w�@[�>+P�l�B`���/�(i"+�*=����p�'T���h����/�U�bmłBܱ�*��ߠ���h�a{Q#��a���vOߵ�)=|��dׄY��Q^�-e��hA�͚t��t�v�ʇ�GN���&3�N���k�w<��{;f���d��l?�6�F3�+�W�)W��`����y�$Cõ�g�n�����1��;��n��}��e�1�z��>-�6bY׻}7��V��1��;ff�c�(��,�3�ԕB���j�mEf��
���fs�Y������Rj1�;k��g[׹���:����� �r춣��1#ø��<-!ޮuў�M���z��V`����כz^�[ �Ɔ��J��C0[��=(�TxP|H�P���Y=7� }%���uH�9[ē��B`T�OZ)�z;�lr���g�L���,|�r�l��(�L*%-&�����/v�{/̳mq����gA�ha\+L��X]Ow�Kß�9t��C��)��b�����G-n��6�<46��!5��(�}�0�.�s�`���� �z�r�~�@%ԛH*BF�[<K�^�	���!U.ZRؐ�aH�:���r�g�%\�O!�+�B�zfk4���P��j\ɪPm��7օ�UFHF{�NO� Q�����з>-�S����0_�e�b��o�w��+�B�J���e�G�85�U㵖�j��V�GD����+uH���yH�YAM�(�ĩ�D=W�GmȊ�łzO��T#�U.Q!,��A��]0�&I��H|��Lay oWp�(��P��C*�:��?c���7��;z$�#>o��ƞΟ��Q�PM�[�p :rsQ�8��?ݎs����9;����j������{,Ԏ&F�P<�=/H�X� s4�-%�Z#!߾����˘�z,-��)kl��pQ��˧T��mi���^��3L<D�8CD=�;t�I.)�����\Ѕ��pR���G��yC�ɥV�%̘�: �����)���n���Ӷ�L�簲�W�j�"��5!�5�L^���ʘ��~x]�jGC:yE� RB&L�44��R�32��z�KI���,��Кi�=����h���##���yT'�#U�w�����
;�C3u �|m�N!�!8aN�}Z��E���S��E� "Π K]b�a��r+����șs��q���8�n��[JӼ�t���̄
�b�e ��/�=r�P	��9f���n�uix�3D�_gxT�+!h'��B�����/fW$��Պ�25��V��S���d�$�L��Y��$�08 ([P.������r�՞Rb7�A���l6a���pGAF�J��+Hlv���+�Q�.�9͈�,$�?�E
�������X�ef<1@kE��h�C��}�&�����{��޺�疈H��A���-��V�\	L�aº]��h� ��,6�Z�r��e������I2G��C��rj'���tr>�]�¢�mg�.�v�x��x��'��4����������)q=����
t��50sv��0w�Ĉ�����!�m�d6��y������Gv�gNA��^ksN]�U=aYj�4HJ�lf�qtǦl� ?�moD-�X���-/+4�)���1l��R%C��-�M���S��7��u���
> ��ȕ[O��+��=�!jo���U6|��w1� ��L1sI��Of*�[hH.�ۤ�v4�ʟ8h�N��fQ����:�ܷpB���H��۝C�U�9i�n.DƂ�]��%�t���x����Cȳ�U��c�i�w�˙�q����)�j�>:qO kg@�t
���r��u\��!��x�r^��Q�!e6�u�5�+����H&,�&�p��R��!"8�.�Y�,UE��G	������#�;��Z�f���߉�g78}��Rҁ���P�bD�-G�K�� ��J�.�NM鶬�:��m �A�Q�7\��B��r�:�;ݨ$�LW����؟����YH����,^����ӎz�x�^�~
�s���~7'�o�r�1b�.��&�Ҿ#+8��]��F�-�����\�H~ ���O��2��$5���4;$/���k������-�8E{�T����O-`������H��w�q��{F~�#��b�6�`�%oᄗ�k��~>��%I�Q��D�"�נ����R�p����S��?Ȇ�̈́q�1s���љ�T���0�w0�١#6ϛJ�ѡ��𗕘G*6��6��ӜW\��6����>��Q����� ��I��v�o-��';����w�OKW���]����/��½�*(��"��S�Ո���E�a��l�E��ν�+"Λ����j�?��S�.�R�	6����8d�kK�d���5�����,��@7��/S��9(�C��mI
�0>�(5d#}U�K6�k��y�%�ҳ����	�� �؃�D���D����yop�])j<�B���4��H#�ک���Lm���ή�ƒ!ŗ���#�l���le6h'xbd	X2��c�i�vW
J�����+-�I����m>>�`�NL@�ӣ{��<�n�)�H���M��%�yt�D�}-��$��5�Ƨ�h�g���fE
V��{�6�/��Q�(�C �4	Bf���|������5붧J4��K��>�[65\bx�UCP��b��F����.�^��"63�(m�d7lg�ָ�����DYMs(�#�oh��#��ÅYhP�������+��Pe�*q�u3	ӉN�)<n��x���	��E�t�LG�>q^Q�~���,�3~����� c�^�N�O���'�x���K�zb��8"�����A�Rɻ&�&0��8^j���0ҥ�{}��rf((���G��#������q��z8B?�T3p*����d��׍~v�JQ23�1I���~m"�R*0�5���d!T�mV��� �`hnN$V�����ҏ�yzI��?	պ��M9Q�e���YU����4�����in_�*��<�p��;�z4:'����-�8�U��C���7�]�bU$���G0�m�n���S\f[�9<t�ǔ�Sp�Ny<M�C��]���ԫaY��7�-�y.� uS�f6�z1{�߸�0LU9,�j��'���C��������*hX�h���(e�ί���&N�K�^��V��L�h��)�k��s�o���D�N�ÝX7C
��}�l��n�d��{��&����S�wE�G!��d���ǒ�Mm�G���i� i9�>�|
���l:���Fg�IS0�jr�K��5\��ݞ����J�f�q=�y}ܮv?Td�?�zW�,�ʨ���u?�	�O��U�M5���	��z ʋ� �m�l�D�M��R�zϩ~>�a�kd�����@Tۗ\�עtϸ|td�����p�d���B��r�������S|kߝL�X���a�R���J,!`�p����`7Υ�D��8��2����]������ց�m4�&H�H�?6 h�욟����%ѓ�$o����Xg��iw�I�{T�8or-;:@͔��>��wj�-��@H�m�O�4i׷2Y�� 8���,��5�ό��b��ܕ�VX�q��@RvR�:�_�?2�FM#�'��Եu��Q�r�� �e5m�k��g;ɖx2�.L�S�J=$�Re�96Gm�^��R�G�va�h�t�����
��^ƶ�wI8�McHDb|A?fG)x^�Sz��yIg�)�o�L�ޔ^UE��܃�n���K��(Zʖ�2./�k��3F0Goo��j$�׍��<��z;�]i8ܦ�U�@�,�=n����C��R���o&����WX�4h�bL�ϙ��Җ;B,3EʘY^A=��:ǜ]�ۆ�[H���f�п2Z��N��Ɇ�tI�e6�-K��V��F8��ܜph�����$m��D)(�Z�6gK�t�w/��p���X7LA�x9������\�����᥍*��)M®�4zC��\��z�o3�����8�.�i��v>ߩ� p�ǀf���rCS?�M�#����̷W)���`B���Iϱ��a�w�`}���9O�eVb��zQ��^5a��Yx>���v=��s
�oab�ѡ��5ϵ@����F>�u�n��_�*��#V�@;��R ��z�BDzd�2�����ߚ
�M��j�^I��k��%g����E��6_��tf5�ut��)�j���oaվr/�1F���]�&\�-�����?�gn�
_�����	x�ug+��Oz��ť*�жG���K�2�쭐��+����X�p�E���O���7��#��x����Q�+��Z��[D^թ�/�sA��yդ8�Y�p���Z�.�D0]~ �芁��;A�U�MIӛY�X��j`{3���FX�����,p6��&�a��_�#瑑��d���*ي4oA��X�>O�����l�VhF��q�f��*Zgf{5L�h�W!��}	t����2������7�#(����_�7��l�1��rί]����g�b�1�[B���	�w�2�3oBo���/pR�bT���9��7��vF���߲��ԯ+Y��])�?��_�Ã8��H��nO|)b���ͥub�_>�1���/���EҬ#<���LD~좩�H����	"�Q�)ţ!��"����.��� e����Xk��1��>��;�="���IL�L��S���K�|j�1���P�ebÅ;�G�E�?jȞ�#gΑ�VM8�q�[�Mg� �o�~N�#�Y/����e>,Қ��5_;���saĠCI7�Q�:��4�z�D.� �d^�5ϥ�W'd��m~c��+�n�vaS���܂̧���O�pV���*�|���Cj��0����6ã��m!{AްȀ. g�ПO��)�^ځ�P�r����fs��K�Y�.�������CȈ�6�MjB6���PGI�(K��%Q�Q��/Iњ��H�V˄�+$��<ai�Z�ۯ�-�9}�z��~��Eu5b�VGp1������b�e��V��Ⱦ��=U�Y�S$`BP�\��̬��}��3�O���mElםN�Uǅ_|��T���W�C�ƶ�J2�w��&���ق`M42_�j����_lO���y��V2�-#�Б�6�_��ue�?&�%��Z�����`��io��ѿɺ�.%��� $�9	;a�M���,/����U�#���0��k��?�� ��q�o|{�hq;��z)�'��5���?毠��(�����{�}ŻxQcW� ��e�zvq�a��/d�a?��@k�LeI��%>јf��`T�'��!� �/)���3FU[�-���	��W�#>r���rߗ���'��YB���~ ��ص�`�� �W
��-G7��L�U��~�9-)m�7����=gS��V}�b���N�P�_(/őS��$Y|�x�`2w~
��CT!��߲+ZX�����c��O�����#(�����.��k��Q�b�z��5<�d�iz����i����O-�
.|)����Tbu{�H��J���;u�=dX�΁Y�k	�ە?7��S�`A�E�aˮ�N� �6�\�l��
�=�#��P�,Ly�����lT{����BT�����Dm�	X�b;��Z�_}�@5�`��IU۴��{硉 ,���.Sw�sp��n��7cj��@�B���~�x��wA���DXap,|Au�cG�Zo�ey�yq#���!lG��"�i��Z���:	���~��<<��0f##�4��^�\	����+��~�ږY��9�ݢ�a�J�/�4����\f,h2O\7�`��8�T,����U�z����<8$�����7��9�^	G�r;�V�1�.q�ϖRQ��$���!�n�i#XZ�(��y-ܩ;�{�o�S?��)����.Xa��؀l��_�=y��eg��_�f��(�_,_&у�ɍ���sHb��w�{RLJ	�e���S��0��^�[ڶ��_�y����q��x��6!�2X_�i������ܾ��nKd��&��P�t&���QJ5�!W=��s�I���=S^��
5�ʥ�a��lkz��hy��6:�j=����#ML>4�u�=�!"ƶ�]��S�^���T�C���
�ɒ[6����/dquk���f���T ��8�}��"��Ȩ5d�NI��q�\�� 9����-VIӈ��Z3N9Y�s�����Q@��6"���C@ro�'<��y�~�� 9Q��������w�W{(��Wc��P�du`Q�=ɞ�^S7-����$�@P�.��6)�����55r<B=ޮ����΁����̅�(�ٕV�;}��9Nq�>�Vc�@�:ջ��Ķ������C\�z��Jrh�'���� A}�g�j�=5��?B�1v��z�@-��8�u�n*�{j萇c؋�4(�(��� ���kܕ�iE)4��z,�p��DGq��^M��� QNG׶z�Ը#�!mZ-$�.0C}��^��=2P��k�	�q#�Z7���ZRt��LsJ�㰨����-�a`|��]R7��Ȩ��Q& Օ�8�́I*�v��V)8���ƍ5�q����ܵ�򅘩�a�cxx:�4A��0�
oKd-0:Xp�7�n%�D�{�$m�u����h�6j8Ipz݆m���?g+�؎}nKA��Z��F��ZN�6K��Y�ݞW��#�[�dGT�!�*@&����5H�2߼n�޳�;�\e��,�74�h�qz���YwDK�*�o�|-A˖}�-�)�-�.�cL7Y�ݯMx@H�l�os��q�
��f)&��C|F{��X�E.���5�ݴ*[���wσ:3�t�M�5�%6��w�B��o{q��D���������%8����π l�������
��1`{����w�w~����E-غA|�1�c�)��քa�A&�e�D����=�߹LL�186����X�޲����d�9��曡YD�)!�3̄j����&Ĵl@�2�C1��^c�J������bV����[@n��!�o�&P0OoB͝R�n5��������$���4#��R�~J���rð��1!	��u|5�zS��N����s��0�X��ϋ�����קt����I��0��tվ���"^��J�����dh��yU�hs�� ��t���s��M`̾؜�rь���`36���i�1��!��ȵ ʻA�Ci��e�u_��2-F� �<��_�6Lꃈ/HRC�]��g#�H�k�� p���_�_Z���p��ۻ����pǋ� ��Z3xe;���>/�l'�v&�i��i�
��2�>�4�1�$��f�pYf��\Wu9(��L�6�)D�K$B�5���B�g�˝C$M���]��\��>kgS-Q�2%Es�)�8䟆bwD�~M��;�>�M���V��_~����6�o�R��HF��gq-u=J)�&3%ƩVW2|�fi�����m� �9KJET��tG�*#��`˄2���c��'�k��ܤ��(������A�������M]�&��Xc"��X%Ly��g�$�<�=!������E} ��Qr6:)XY�ӸW�%N���]z�9�M��������L,���J;�3?ɢ�W�_�/ Bճ`�dv���K��6E���sN���Et�i���.$\��~�XvB*�X6x릁��1}��@�"4��,�啑'���%�A���C��ӈ�����@\���Y<�0ބ��hȖR�P=șɜ,�Q�-�o���n�S�GOM����)��Q �o�LJ�q��������+3��i\����o�a��P�v�H�����'�xM^��5x�ؑ,3h����I���"֒��R���F�p�}��a�ӄ�]�ZM�{9y���Λ� ��^=��"y�*��_�2�#��Dռ.7��L��>S�����:ь�����{�O0hg�9���9�+�
B�X�Z"]~l�,N�h+����;Д�k�q�˾�f���Nƾ�v"��gP�p�A�(8��;�3��n2p�SP���T���0���{˻�^���ٻ����u�d��;�Sq/��oR����R|��<�L3�A�x���-�zh���
/�tAe>�W����d��=��o�Z�w�x�m8���6�&����$�����NY���r*<��mULe�j�e4)�p�(g�tȣ��I(��D�}��s��Mͫ���7i����&�}�_H�\��}��*�(/�hli?�iY�FB&���V+O�~	�Q��I[����r�������ܚ�\�:��}�e{�yfo�3���d"{�\�W��C��]�p��Ycrb���f��� �m�.|b�����߅c�?O��eD�_��a�]�J��~[:�#���a���`��D�������D�Ԓ�;�SeJ�ξ*��X�o��1���e-kgu+���F����Ǭ�7ӳ��>�{��<?�:EPe�g���Gy�.)+wΔ�F՝��>6�>t{�v�uȥ�.aƄ\��
؎�����e-�
��:�
�JY���� �P��!�r��hٯ�A�Yz�L}zB����B�Ӌ�ĵ���l��Pjܦ]�@Ņ8[c�X꼉��T\\�,��~��3��Q>�!��[��t�K}~��[��>O4��T��p�B(6��yZ$d��E���h��h@���dW��;�=J���|;���+�%Z���𜓒�w�S�ο��]u��	��h9Y?���%^�.��F�]��K�&�Z�{�;8(Lb+��zBP�Jq��d`'�f��U�R�f��HXw�?^;��T���Z�K��x��CH/��-�d�:P)�3��ʢO�)����z�;�hyj}A��[̊�Z��`=��ބ���O!�C+���p1�Q�_O؊5\	Ӓd� qo����Zj�u�zu���"�e���16�iߺ��u�y=�ԓ�[����7�j������c�ؠGTK����!���pVr���y@d���zy�f��K���C6�>!-��p�(����Ӳ�qz:��Pb�E�f~ t�4�=���?����.8O��\�ʣ�Ϛ>�6e�ù'�����뱦z�H��n<q���H9���̰)p=��P�߲�m �L�$5U����@����	�|��2�Qk۽�G�Q� aʼ$t�xL�x��f*�������x1!h�qC҆3�$?ֱP��f_���t��ד�m	xI�і�g�.�oQ�7�fϼ2=�KòRxlo-*�3|#ir�Ժż��kJ����o��V1�9�űIjdG�R�F��wUPʐ�j��{^�2$R���-�A������!m:������=���F������.~^]m=���.1���� �!��(nL[��v�=��0B)0���) �L�qq5�����s�b{���L���˾bv;�TQ_*r�'|��g'�T�'`mЕd$���h�&o��
��1��q\�Nt���Z�ڳ�-c���D����J7ry���#����U�[#�
*W;|����2���)�O���O��oC��mP���iz�|��y�#�JE�'��J#:*O�p�w��NhUHk���v'�w�V����+k5�4�ņ@5��	
]r�n�?βVb*,���©p1HN��r繻ӈ7L�J�E\���_@p&%��3%�O�7�/ݕK��_��䶪�װ��#d�_�lijC ̓��@c��(�^�j�l����<j� ;g�p:���<�[�����(��]({;�>�*�h�&0�ζ�"Mc&6PN�!����n����h���ӌ�{�a��5I�I4�G��2iZd�J�)%��Yލc1f��U�M�:2�7�F����t�xV���UJ��s��,��`�^�嘟�Eq[}���f���	��{��M���p4#��⵽�4�hYs��8n��7�L�Q�RĎߩY��L�E�����et�gi���
�5��ֽ�ͼ��Շ�D�h�#\��p�QE���;)��Z	t���uq�sM;BZ�5�7gg0�@�a<�m�!Ј0�N����پ~K�v�+�r�O��f� ���s1BH������ӏ9W���,�n@vbz8�	o�r3���=W:�+}�#g�4N�� �x7����|�	ј��pޫcd���޸K��{G��5n�;A��k���D�5w5A#D_0�~���e�:�$h�<5-=��K4����]��2���,w�s��h#<t/�8s	\��%�b�"��2��jX��{ˑ�>� ۵G� �	��M���mMA�����>n[�ƫ��B9�t��=�ֈ��AQ�Y<�Ģ�5�*�������<S�9�o��8K��O)�`u-`�-!�+2l�j��R���k�%��|u(��̏.��rj�,�d��fEKp8�l�"��r���s�,e��?,�� {�G��_%�����>>g��R���l��)��$��C���'9ȋmy���,�TOrm���Wl��wCn��R��MҟWaK������i �5��.'>���R��I�Mʾ3��q8�AOV ����Ȩ��I!��f&�5�n�ڝƔ3l�V/�B��u��s瀢��Us���#>Hr��w��js6Z���ʚ�̒�%:�n��_ļ�E+���Dz��U��� ������j�o�q���o����y�hqo03pbcS���ՁCh�� �]q�B	�M�
�]�ε6|=K!���t1�c���a�4��a:Q�kcB@�-(���}b��5�C��Ie���BM&-��{:$�4��*i�D��C�Z��=�@S�G��
o�T���1Vb��b�����P{�q�>2��E� �@s>�i�/f�p5i�ck�K�f��`�7̭������̊U3��$aI�K����5�\�"�ߵ�mM$c��QY-��u�3x��χ������oҜtZ*�	@��ܿ@�S��[s�]���;g���B�}�7E2�C���13$
�
��/I���`��f����.a`T�#������<&�x�z�KG��T,��B=k��}!�&�y'�ZH������˗
�� ׆�̜XQw�}׀[���Nj�J�� V�~�{�mB�C�Q�
'tw@��	��}x|e2��OG�vG��Mrh�=��5����f�vM�:� ��	q/��'���+~1�*�|� �eЎ���DQb�������^�'�W�X�B����/|�.�
#��@�5��NK���Me`EQ��F����7B-HrQ�m�N2&{Z�=��吏<�Ñ5�!.M���b����b��@�!$zR���KZ�{�����2�H�m�pd��^x����>F��%��5���Σ�q���ٌ0������O�����\.���2�+��hA(�E� �³:d�a�a���쎸3�M�զ��"C�x��񚅫t���֤D9���Ӹ	��~:E���zWG7�pPG6,�6T�k�d��O��rW���Il:�q�~��1~��������:#02�����M7&��M��q�_Ȝ�6va��,��:�8��b(�*���}Iq"�̨g�v�DT
4��L6���g��<rHA[��p����w�鲔�i{U�ӌ���c���[�$�7��,�j�<R�:�K�`��5����t��9y��r ��r���%�.v�UJ[� �M��sU	�,Z�yy�0�jL��Z��3'�ù�����5�v�@�����}��Ѭ���41��i�@Mn�	ڳd�-a���lҍ�ƫ�u�JȂ�X/�و��[�a_�e1�b�f���Ԯ���d� ���õ-�$�<g�=�p��<���3����噘jI
ܚDQ�}p��;�;Z��x]���ѓ՚	��[ju/��=[o���� B.�O�+g)�	�ؤ�o�u�u���E��1ꬵޥ����}\�׉'�$%�9VzE�p�p��IG�4���-͎�0�0�yl��(פNZD]��?�������0$��"��G
�%2�t���
۔ϑ�@��s,Ɏo�,� '|>'��[�����p���;N�iൻ��{$�׆��E)��<kx�XIlX-�jS;�e9dbΤ}#:Q���oE��UK�s�ڷn>���/�u��oD7>�њ#���dE��s��X��sȊs�RW�˹5~P�1L�oF��'��Q����"]3�4�*�ۢ[Ԓ�?{m�i�A�z�#}B�����U�J�G���P�f�d��`�2p���r�XѪHF�)�.�38��Y6����LԈ���+Ȃh�B��a}���>�	��ȶeBٌ,���SI8/��^{m�Ne@\Q� 	��I�v�)���#fs&O�t�i��Tk̟���,�4-FzEq��9���?�S��L4a.L阔3���l�-VUe�<Dԝ�V�ASƒIH���=Ȟ�Ι�o=Ėw!�*��dr���� t=��ec݇mR�8l�6�,3��������}���.�荣����~���^$�;0��`��~���[C[�f�{ȡ o�%���a
 ��K�xv�
��c�ad�����.Q�"�_������a?�E��lg}�:]1�����)�gg���{���*@�`:�+u.M���p��GcYQnkX��J��܊<�%�y��4W~�����s�m̯��#���G��l�56�l�8�bܔ ���TT}�&�"hT{��|!��(�o�Oj��6�ON]�XtW����6�"Y�����V��#��f/��4��>n7qZ��|)�tt�uߌ����5c�[��)�$4rw�s���I͑�7AľdoAE�E��R'b�S��S������c�/>R��q�;����㩅+��
O�\?x4@rks(�tI���ϔ���և�*y���+7��{75����I�wX'ٰ.�t[��/�6_�J���ţ�X#����$!�p�e�DO���@	�~��X*����Jc�ܔ��\n�K,���"f����m��M8��1��]��-��(C��6]9oҊn�	T�D�en"�<?�c�H/���W�A�/��h,&Y[R����c`��qah�0������6E�}L��c�*A�C�׮@�;��f�����US���Lõ~m|k5w=�%iu�F��[�u�n+�R�����Ƹ���J6�I#Y��`pm��3��I���Fպ�e5��a��a0fC�0b�)��OCYB��⌖��!��!��	��3�X}��&�5RÂ<d�%!�m\�i�AD�m쇎w��F6����[#(�݈џ�\;���p�p�;D�y���}&���q�O�J'h!�:����DX��j�R:`��6��1s1��L�VT)/���Fj)"(�B,�#��Y��da�u�J�5�*�z}��l��D'���9p/�h�TF�mN=���L�}��i�zM��bT=o�/.QBD�8L9��7��m��USNSH������!Ʃ����
�^��9 �,-����	���ԑ�EN�{dëCW��Q���M���D��H�1b��ҝp�*U��y���A����!����k0>����~6Z`�* �4H�좷b�<*��I.��,xJ�3�҆^M����$Yi�sc|EM"��ؘ�i���+
��nM��b�����'�X>��W�Ἃ.������_U_k&t>�)�5e𣝋�,�Q�9�������zRn�| U�b�r�,\x'�4�d#�9R��fqN��եo�q'����{pa�\�q���=��`�b���z"���al�����$�ݓ�{�9�α���?YH�!��2E��F��B�?f���>�4�pT�El��6H��{	�
ST��f�i,A8T!@�B0�h��?Ja.H�7�����|�&Z^�=?Y岤0���RW��4�E����
���de��
��M�52\���~r1}]��mڲeC��K�]��6���5������mJ������Z��vH��%��]9��,v[�k�;h��� ��'�]����a��Z],ϳ<�q���#_��O|�HQMK���B`XQ�h5�pa=��<F�x�Z����,|��� I^�l��PUݛ���]��~gK��C��n�e%�,"�W��"�1��Y��$���I��w��~`&��B�Vw쥜���1���m�κ��wب���876�������&d�"ob�u>(��޷�on^>�G3��}��Qpj��&��TU�iՍ��>����R4N���s���(�@Υ��S4n-M��؆���̻�%^���p�<D���")1�(`i�B��2�ce�_6u1�>�"�it1�n\~��)ʝ|ӬE̦�E
S	19�*-}ʙ&!�;?�V4�`t��J�2��X�N��J����@��uo]�Q�'����߸�@+�-��s����oj�݉�M�B�NI��3tӿ�7��Qa���ГL+9܅�(���@�5ðm��צ�$��z��}e�j�-ǐ���D��!�=\>s<m��j�&x���*d�H!%s�
�`�����:��Q>?� �n�r[Z����M>�L��G_����W���z��?f� #K�2\��2i��u�}�m�Qޗ��>p�<d ��@!xm�f+�K��4La� ��n.�q2:�{q�� Zќ"> �X�i@c؁�ۯ3����M<�Җg�`��Cn��2O� �%1�M�@��Б{8E���hg�e��������h�W+Oe9Dxc�6� e�)�H�|���S��s�j��v�nn�bZg�-*��g���d[aP_���_O%���Y1Z����/ ��,���}����s	NnȜ�Qm�+ڌ�h�r�@�φ��_�?�6�����Wh:f��ގ��3�r�%�n��!f�R� 	��S�sq��;d�w��f���-#�S�౅��K--<�tw��t%F͇����*:��A1��N�������PKtm��S>v�}�O"�����;|��#MD��e��Tv���E���� u��)n�)�]ی����~��?���
�Y���bds��?�@	�Of���p���I���y��h�����W�`�YϓZ�|�i�[�l�,�;x���� ��S��̒�Ff��3e�?�5yr"���yE������+�t�7n/�Hl��^%�,��a�p>�ZEn���7�O���V׈�U��*���^U����;A� �n��� ~�r���v_�&�.�>ʝ����.k[����%�7n�l�G��nk��b��~�\RK���N2͋hh��S���$�Kʄ������*�UǺeQ3ӑ�d�X놐�N�N�T_�n�_�*����!�d�_΀ΦpA^�Iy�]y3k�������j¬�UkU�Ⲁ��O�B�!w2'�8�}�����w��n6Q��8�~wcfF��5�^i�9���/���KU �������~4�9�}Ϸ�x��՗��hT��U{:x|jPt���H���r�~|�@�-��X"���6>�h}�kWbdŚVsw�(W�6j�Z�6^5��ԅ�dQP����f�ܸ�����.���|~iQ�ZqNB��7��B�hl�!C�@[��ag�@[	 T�!�=B���)D3��Ӗ[��0��H�^�~u��JY4�<>��\]$sz�l���2y�AƱ" nȃP9*A�PG��=أƣ�Һ-��W���G�A<MP+��/���J*Ξ�m˛���$��SRlЖ2y(�T���>�6���-I�'��h�Pu�����0`��	v�f|��3���s�,�C�.�nz��(#����#�W=̀���R�<�mk���>�W	�n,����A���뙿 cg�k���r/3�JݶH�A�?{_�rp��.����c[�ԕҨz"z�e��$��bHQ���}'�mDZr��G&�>јϸX����5[���A�ςSj�@�9�Ͱ�w�ڹ�+�!*�ڤ\��b�Fj���v���FB�9������+ ���d���^�}�Xlj�	� �>zӌ%"U@��I̬^iMe� 8�R�>��7<���1�[�!l<K�]�W�6w�$ӌ�u��A"&V�oR���4���~4�<��
�| )�Z:9G(�AK�b�S@M�j)�"'E��*p�Ni���c��]�hgS���r���4�Z�g��$�G_U9 �2�,˜��i�Gdb����52���y-+��u�4�3S�����}R����ݚڂ
Þ �C��#�>q�h���ё����2�h�GͲU���7��Z�N�Ύ8�3���,X@�u��8V(�����ϸ��X�p�_  ia��S=�=��EV*d#Vy�CI[���" �g�,�ï�\s?�z�hn���4�2�+����
wt�]�gX`O�r���R/����fh���{xeG�_��<t�b�tVY)��՟뺳�jU��_��b��
�/5G&K���A��2�P��)�)0	פ-uP�8��D!�4��4�����	۷6�6���Gd��������_�ύ�̈�����ޢ�,ٷD�nj��͹��� �Km�R��y�:�tc5rTf�+o���e�}� `�`#�;H� �D�HɄ���tLD+����
P��%��(�:B�8������������@j��%�/<��CQ���~Yx����D:/d�Z�����(��^�`��tX���	��)E���1����W�h\�8�h�7�>94����"s��F$��i��~�(�&+�pixW�:��ca'�/Pp����� ��ma�dI�W��|����2�,��v�,�~H���za�q2�fo'�S�4������75�N���XQ��!���8c*�C͕ػiU��5Y�
�ׂZ>h��&;�ȹ]H�� �.ѡ�:z�e�m��}�>��=qnBLP���K�l�Q�v�|#LǊ�� 2�B]�X��PT�A��t�2�53�U���C��Y�Zj>w�֠�,T)D�
FŕS�f�����8���5��m�ι)�H���c�NK+ �*@���H��5T� �r;����p�`���~%%�
�k㤔���l�*~C��迵�����]d��Ѐ����ը|;�gPLr�?� ��;o� �D<F��3t���OR��h��	�:������Ʋ�À���]���|�Tqj�+��ܖz8���<u�\QvX�s���܎�-}��N���L��r ����}�o���<agO39{J����x{�>G�.,+��5�1qQh[r`�L~�FƇ��k���A��r�cx��������~�;��ƇG�\�:org��8Q����"u��b�f;c����d<Cq������=W+���������0��5� �]>�-�kt��L(�8&n<��R1����Q��e*��Z)�S.�$g�k���":VA�T��h��ᗖ-}�K���߯=q貈 ����;�7�9��b� ���_�fu�U[h��AV���NO?9ND�3�澕e<�ܥ�ʌ��`,��4H�<��3PNK�m~�L�(|��n���(l������dpA���{�M+a�D;��$���u�=�4H�	��$&�1!|��f뛄} �@�������o3X�=����B��������tJ�UN��m�G��T���b+�ra�7�_��,���t�+�)|��w�N�z�"������r��@���n�������O �T���#�忡4J�6���4p�8�K��D�U>�V;N�$�De���5B��u�B�� |`����Fq����h&C *����w�=
��Q��2W�kѾ��nb�Z��1k��GK�"�TRhA� '���~N�O��]��غ#A#wZC��rq��l#:ڼ���x�k��L'7���M�P���s�'��|nce��lg~��W7;Y{`���Qg<�>g���R��F������FPmsյ3�vl�P��Bn�!_���y4���Tb���t?�~�`
�V�Ǒ�gg^0�Pn�~�j�-{9�$fHN�.���k"ۙFZ��K��kP�JQ}P>Y�X�W�ȴ�#G�?���>j �>e��&H��i��n�V�?�X����;r����S���bJY�אxg��H��0�����ϻP�G/�UD����r�����x�����ϳ�6�=�w�Vp�pm \ĪJ�ʣ�`B$��3~U��m�o��&~!���;���Ő����6E9�L�� ���2ޯݙ�P���G^&�=�Em
�H���_\:�^j�{:�(��Q�Y#d���<���-�R�i9��8jO\xbS��alu��o"A����	<5���F��〫�rh���}E��@7Vp�w#��y��h^�r [��n�J ~�YO7�����&]�`n�Ć��R��E3Iz��ϥ#���rb��
��]t<s�=9߆���n8�#������"u������4U�$�k岨(�1�S����*���igf?�g0�TDT����;���}	Z�9��PN�GN���&f�R�b��3��x}V9j�p��B�&kY�;U��b���9z>�	��؎N�L"9p��.�X�F�:�.2��U5�/���Q;�+%8��`^th2nv�3_�Ը2S�L��'o��!<��H�k{�F(��̄�& Z+d_3"���n��~�ξ�+W؛CZ��Ked]�xU�5S�-�>��7����\
�X6u<����
�]{A�Kx~y��O�EْF��#g�^�Y]�w�n�㲽,�Z�<M�����hd��b��^u}Y���t�]�������݋0�]���[%� ������떾��fg4�s�Z�ۥ@ �[���2���Y��������
�}P�[Qiڎ;��e��
���;O�K�@�j]P����z�,G�=�Z���{p������V�x����I��]�b<�/�d8$��2X�d�TWNw�w�@��7��g�K��m�迲
8-P��-�@VN����a����"�/�����4��ȍ�AD;�k��(��M��B��[C�d�lp2
_\��(5W�_o��H8�yM�r�Bu���G�5������{�w<e��q���; 6lRə�Wy�<Ja�Ǝ��_�Lv��@Tg�Qvid������)�F���Y�w�H ���Fo[f�6��_>K �BR�<f��&C��g��7�%�P�
��Y���;-ڊ�y�1 !LA�Z��?1�Ӏo���R����(����SA>J�1p&@HP�nٙ�u,pq�%m9�/�X��FU��p�ٯ��޳�ܷ�c���ud�O�� P;2�`?��k��@���gd�iV�1.�.�ӈI��P�HM����9u����Y���Q�<��_��-D[��Aj�q���̆u��x!�}��Q��^��vη�ތO��-|����;۱yR���oH�5�nj$+�ER�=�]]�}�6��GoD?Jy@��ϳ�;�
�$�{5��N]���u���PvA���mz�w�c�O�۹�o�t��4��<���~:���R��^�j�L�K@��m63h�O�_T]��������ԽR��B���%\�(ۓ���ڠ����㎛1C���9��`1)�U�8$f�<G)�4�ld��_dȇ`�Q{hЇ�8�!�Z�*Pi	P��2�����Q��*�yM�n���{����C�D�C����5�8�;��a�Z��(�A��~�g���Y�ڜӯ��ӗ�{|��c���g�M��7�a���OW��.���4�b[�ҚWqj`:��8$���$a��m���,�Pc_4b$v��Z��{I�sm��N��	�a��#;=���mZ�Ad�_ir����Yf����2�\�xkB�"�����r�V7$j�65���=0G�?��>��J�z��,�oV��z�w�֥L����A.m��Y5�4��W4���	����0aags�4B�e�`hd�n�}b�ɞ6߮��6t�6�k*��e�>�d�c�}l�$#b��&?��T��c�.C��8�}�������#b��Vl�褜�
������rf�&����)	)�sPɣ
7�T��ݿ�2}����Ø�|Yi�L/# �UF�#��x�Q�V���W�<�������d5+d�7P�oA��_�/�m"W����i����^���7�t��#���35�.F�`��5d9�V�m�9c+�~y@�-����a��F�f�ƪl �v��ST�^�t���,w�y�e�:0e�TP�t�ލ�k�ӏAA|��I� ��"3�@3���s@ƜϘ�p�s�+7��T�k�lx�J��uw��]0�.���2Ͳr	�Y�(q��R6���]�N���,G�.�@6����AbG��G��ާ�i
+�0&8L��s �$�Ѳ�Ҫ0��q�K��y5L>����H��`vV#Y,C9FWQϵ�v�i�*#+�<y[�=d٭�i�L���-�pf��&0��g���Ϲ�#L��à��m<�q�A�d��*�F:���
�T�tm�v�^�K�����f�_)�fOn\���h9���)2����P�t�@��:#e9���{Gð^y�I#��M��iyX�1��|ו0A$� ��R�����^v��n�
�}���DѢ�%�R9s$�ԗ�NŎ;�=k�^�[����@�Eĩ�C;��:4G/��ξ�ټ��Y���J����	����J
Ů��C��H q%CމO��Z��D��F���~_|����M����n����u�[߸-�� ֛a��ޯ����<����Ǿd���aqH���`�F��Y!�1�j�X-	([���°$~�pë��{m0�~啠+��ȭ��M�(	�Ͻ���"��bz�2q��1��gD|#�Q�;3�M���3kؗ�(*Y��:7��H�[TQg�BS�y*�ᢲkl��l����_Z#rt�1��L΋��bXd4q�YH0�v��6?D���o���u!��w��9���Z;�z�o�y �Ϊ�GR�a��</�'V^:������o��^������l~�e�ؔZ���M~mEa�2p7�D�Y��?���
����n_�LPg:�i����߮��:+l!�	�!ҵ�"Yodl��|,��0*?�?�,���eW��7��Q@�d{�\ݪ�����c��d/0h�"�5a��!�龭��-�jV�<��pI�;���i{��?�㒝������z�K rs�t���ݭjM��Ey��s�Y$��Bfg��>��q.��fgv��xߑ��XW�;����\<	�?-��u�ViB����-��o1��lOU5^��xü����ZHK:�ȯG��H�.�h��(�j|�fKC�8��+;�x�ǐ����M0$���1��e��Al�ǫv�P�t�_T�p���j<�jc�F� ۖ��8����N�0�C��+()���9=���&� �m�בB����x_��d�O{�2z����mZ�$Pa0xma�[/q_�@��c/��`@��r�+�R��}�>���Te��	G����{W�9��U,��Q���iz�s��|�F��c^����G���Ve4�s'`���;'�'<�y0/�<�DށJ�p$|��K��ƊH���;���ݓ�i�}���\Hloi�x�5���=��}V#���d"I�Y��y�pm���Yф�؀�k��*�F}�VV���$�8q��Y<鵥�	�{�������G�
��̢���6��UO�Z�����?\{nA����\���s�@[�v
��xt)�a��h��d�m�^�9jz�Ȁ�]'\gVF�-C�>Zœ!��!A�n&Qg}��8����A=i���/��F+Gz�`:}+\�H6rP.}r�D��LP�"���ﯦ�s;Y�8�5�ԛ��5��,���a� ĭ=��`�QLA(�1���Dfs]������>C��!!X�ӫ3���B[*-c1�gO����o�1뒰����k7<Q����ͱ� �=�,��/l��h04C�y�6�n���#�a.CW�.���muf�b��I�)��?2���9��9�\��գR_6�bo�b~.P�sR��1j��K7G��Ԩ{3��N�zp���H=�q�ײ�����z�mk=�z��s+4&Hw�Y�~�?�rPH���a��Q���y�����5��w�T�_�vA��ܼ�*�&`iHq�|*�.���E&>����J|��
�o��r}b�p�:�[�hR\5�s��+l7E�l֧�17�����"c�yE���.a�ٕŁρ�}���g��#m�Q��k�ȓ za`I��"v�� 5A'ܕb��ZDP%q�������oV�J�@�{۟���b�0�vX�A�F6ߊ���q��f�/j�²R\��(E�䜭�t��O�>kxھI�ɶ�>���˭Zs/ɫٷ��|��P��S;0�c��ϳ�˥~�}߰YN�s��jb�_�H�/:�z˖�f��6\�t�|e���2�Nt�v��9�]�!�4�m�n������e�z�mF%�{��{��A�91�rW���1nSr1��o���T4䕄_3���z���?'u�;����Ƅc��H���*m�+&	�ж$�8�ls)W�t'�)A�̥0��7����;-�����J77{����Uy��F��x�}�]g���l��h�_��h�
K���*Sx�'N���=��g��KO�c�c�[�h`�j��1G��2�v��Y6sm�?�H��_�G�%!�!kXKt|����� >��i}B����#�=�c�Ӎ�z扻�Q�GP��gŢΫ͔�^�u��	u�Dh�����G=�+�#/��$!���r��TQ��Q�{<�mܽ���ߚފ����;{�`�آP�eA��Asqb�`��X@<�y����/�[�c^�pp�� �'������/��'tt��٠�C�d����@�d�1ХI[`S�a�m5k;��|y=�=����th��@ƠJ�Z���	�Oη�v��g�r����Ϥ韇o�c)
�ͧny�T}� �M�br҇3�"��b�7��$ �Ǘ\�̩2��A�w�,�����R? ��5��?���Ko�=_����Q�P����Df�~�\p�%ޔ��݄����@�>��8��r�����@�ƖB�I��������h����SْĲ�wKK�A6~�3�7�/\��5bACr�%�ܕ���ܸ}ԸE��nT8���ިhb�\�ێ�F�	aǓs�rH�<{c���l��i��b�H&o2>��x��FX��s��#�������:��,C�n�h7a�fpl�,����~�N9qKD�-��<�3�m6Cg'E�p�,����P!�ﭱ⢙�#��'� ���7����R?X���V�;a��U��VP���cjX���;�|��=���ɂ̕b�ʋ�@ �L��_Ʉ���^��ӈXM����^����t����#L7@d>���i��'�lŽT��*���8�~7#��"�S�}�,F���=:����~^0�"�&X�Fa�ڤ-�sŮ8c*v��m���"'���C�M@G|O���`����F��n�p���[9Go�t�{���	8�}�q!#p���38HS�P��KBV*�03�J��v)���hn?~���r����!�LP��k�G�C %P��!	m��)�:E��=x����ET/����"�wS'����A��Q���,7��>F��UB�~�l�����G�Y�g��a4�o@"���ax|��/�:y�0��������t��I��6��x0�6�p��v=A88j������^$�FK��ߡgʪ���||J}��y��[�
�SE�D�U�z�  �����v�<?��ϖM��)��C�(�U[�2r��IrN��	A�^f�5�Q��[�l��g��~�L�(�\���RdMm��I6g�����P4�wsi�j��e-��N��ߞF@*2&���tײ�'����k� ���w�f�>�,��9a��k(����ޓ|�i�rz�'fdX.u�O�̓��:1��ve~��]���]�O��*�CvJliQ��Rm�G�q��~[�\�D��Q�Ɛl��ܜ�P�t�}&ӊ�X7tz}d�لh���zi�P�u�vPj��d�k��0X�(D-P��ՍB<�ks�ר�u�m���F�{
2�����ڃf67wΗ(Р�a&�����o!�<:,�%��wFr�B,�
��D������=�giOm���m�*��{��FaO`2`g��f�TZ|������dq�i�� +���-���Kz�G �?�Y�.�K+����W��ێ<J�4����
�#b�{�'� �{�ؼが�.��%��|i#s����ʿcw�T��I#���5zkqZ�G�`���PW����BJ=�9��D;.��TVr��[E�h��Z��7G��&�S�<�G�ĵu�`���\|�N��Ab�p@�!B�zAx�(k��HSN�=�R�7�Q���b�,��O��_�n$�r�GS�.�x�9�;G��%6M�Q"�,�� Gb�I�KC���[�d��,���X\��G�uxAv������c	ī��n��tOՈ�i(ف#�9v���g�ğM���������o{���j�*�f�G��=�oh�G��v%=>�J%�1��,�'����"��m�J���"a�-���<9;/t����8�[�d��eXs¦�J���ʜfi
뙻B/�W6��-����ǿj?-�##�MCm�sez�0)���C�2��Ջ�bD�ׁ�xXb $\�<�AŖ'({P#��Z�&�&6�[�[R��"H�k��S�N�t!��4�ఽ���U��:���#K��Tfͫ�iz�
�1WK��P[�U����	7(�c��SK�����)���9o^��$$�^�,�
<��d��m� q���ʂ��Ih�X��� ��.u���2��3!�`�4��TT�WX��W�= 9��p��Rޅe�@�~)_"םXP_[�N
o1ۣ������G���
�U���͞��c��?W�c\���Fn�!�� ��uh�vM��������	���!8�F��Q�8ZH.ynd�to��M]��p���(��T}�8��:Sܿ*Ҵ.�y��X��p��jk�h���Em���<OC,�w#��D����6����}�a��%I�$�_YU�������\����f�M����m;��'h}���딴Uۄ��q�"��~�"��4H�:�����s7��ٙV��#�o@��xK+��y6�n��9��Bha{bs���&"St�B�0��#�eI��)dl�.�ߵ"�t��R��Yʹd�x�mQ:z�Q����=��(�V8%�&f�>� �|s�P��
��������,4��gA�Q�|Up��6L��ݎ��v(�}��g��p�� y�}Epj�c!���K�a��Ty�w~����BM�M(��^_J���X�tZ���vf��Eǳt�o���i�f7"���VYȯ�s�S^�W��zq�'{���~���@#^mi|��T"#(~)�gz�[?Uq��xI��a��C]w�VI%�c���`V;���5{�`�=��[������%�����*�:�wC���Z�\�~��������}MS�_� ��5���K����xq�H9i+Fl`ծ�%{֍U;1�'.+�ll��Q0N����W�>�qp���x��+H 4��%3�ka�jd��W�s�����4	�7�eb�m?9����1�3>�R^*A�J�E^�s�D��o�x&��I������*�8������͟ˬz�xL/��ќ�b"���x��D�ܢ/Қ��3�����s����q�k�]�!ᤠ����]�������b�T����7hn�/�N2K�E��q-�l �Vjr��(�"�J7��4+r	���.b~�Z�R cM�bH#�Rc���V���VՋQ�U`YK�f�V���I�5U�[Ɠ����a�!p�����D`��'�(Χ��,Ftz3�(I�	"dLه<��Z�(�)�+H�0@,�Pd��X��\˛�R��{`&O/߱ZG��
R|�6�}�����{<� ���tAE�9Ur��-���">k�E�h�#ޯ ��+n*�~�qh��(�@<���m��D�R��l`��.��OD�8�,��w�DG�;�t"5�)�܃���@�uq�SV����ӢW�ߍ�ȶ��ì��2̿W��F}���h��ӡi�����v�s?�8���Vr/���YH���[_!k��s�vpk<��Wb�t�K�Ad"Z�2��gxo:Z��3��o��l=��O3 �-h�=ށ��~�~'!���$�.�~�-����|���ë٠���)8�-;yKÖ����27Ba��H,�ق7�#�9G�Q�[;�;��������xY˷�ݯ�nQݞl`�@:<z(s'�gw�����gqX6�k��c��[�)GF�j�G^�(]h�#��z�`ꛨ 89Åw�s�c�U��[�LK�)n�q|�z�����̲�o�~��9�ږP\��Go؄��%ɰ�l`�0��R͍�gTB]	�oi���iA��&N(����C���Z�V��<���0	�A�g�PF���V>	�L����P6�6�U�5�M�F�T�H��@�ZFO���F�u/�Q�o;��~� �/�HԶΤl�{	��5��p ����B��.B���O
�����$r��	v�"&xmap��g-���n����r2O�-.�[m���Oi�E0�:w@;��(�O�
��J3�k�ˡ���K�jY�}�m �n�^�vlj�}9oৄ��q�)�<�!i�U�!R��J�Zy�Z�v�w�W��n:k�}�#�z�1W�H��}e=�ЌLQ�J��o���ȭDd$&7�Q�%����QOz6|쿪/m�ܨ&��X� 9���*Q?)-�b�c�:[��d�%_�����A��#���r�H���E5l5 1��%l�qW�q��t��Okt��tF��E�Kc{�ɽ9��ׄ(B��&���	eB���W Ͳ�q���3�X����Ȓ9m˧�2K�<��Y}}�G�.����?f�?6*��=�p�k�b�jp�U0֥l3���L�"Jq�JMfz��~����c��d��m	���u��}da�S9�a�ۛ+1�A��Ќ�H�"�J%�g)��u���\!��ܐ�S�fI���ܟ�"�����锛�9n�_�i�R����|L �4y��2�skr�6~9��D;H���պ&��@���`k�ɭ�c�G�4�?l+�B�r ��c�.�j3AEo�4�x|��siKB�[�1�_��#�Ma�U�F���G������<:'E�fi��RY��@�R�=᧼���լt��X�����A��K���{���Lq��<�w����or0C!��. C��(^lP�]f��5�� ZY�tE]��r�J�9e
�|@�z�1�u�������l�2���v`�a��De��	<U�m^?���}�n�e�<�f��IA�3U��9~��nŤ�L�i-���|�3��y��qu�a�ڙّ�r�t�M9�}�� �X�i�������#���ѯ�������19���*�>�\�1|���׸|�L�-�@}��D�M��>Ky���K���G����x-���c������tB"TO`Z��}�ar�6��	���۹|������۲R���;�z��{0����lk��?
��2ȶ�0JE\rbÖ��h	��1�5��N���M��۠^�~�*�/�oo�����	����hy��Y�ݳ��M]s�(F�c��=W���9R;��g�i[���]������^6^����to; !Ϧ����K W����-YK��J� ��
*���n)�1��.� נ��j;�9�x�xӯ*�`�|�/�F-�$�1��e�F�͋�%���:�3����:f��	��&��b�Ǣ�2��}/����!O�N�h	��Eu�]�Š����Z��!�xC������Xꇑ���a�_,�i&CӑxVX	7;�ڽ���Qn�!@D#�Dwd�CsId����}ڱp:��b�
k�N�QE�L�q�huTk+��O|�S*}i�¨�qb,�w��$e�$w=�t�0�bh�_>�׷z�5��rr�V׳���G���.T����NT4D�&1p�Z�DVh�\ג�]%:�\k�W�ƽ�\πM�÷0��(3��֗�4��<_�i�0�������*�1�\A���<�!�35�����Ǝ�@6���q$��3be�G�] JzPO�]$vB�x9ԨPb�C���˺S��eL�� �E�5_���-ξ�Ua��ߘb�|�����N�w��F+&6T�*��G���T���v(��;6h!�-�$�hN"�3P��Mz��0��@Ag�L�w���u=���r�ى8el��	sN��y&���E�e8 ���7�E�xQlOp�_�%�L�d��{ۯ~�h���dS�r%�b. ���k��y���Q��K��`�.���8�f���ԉs�1��,�������Z�T��M�N2OF@�)������\r�@�R��4�uwjth]W9�T�kM	�4@v[�I����yף��|�6;�h��/�:M 	�*��R2���?�^f �1�d���)u^ �,��d���1������!��*Bw�T(�NE_���� ��Ī-�T��r0Ke��g�dtm�"�(�]*�l���ҧ��9�CcZB���	Q��9�"rY���f)�O���tEⴧv�qzx�z}m�B;d,���d`q>s'6��������?�c֋j6P���*���q�5�F�|�T֧D�'צq�jTr��b�ٴ�ʧ,��GO�k�uò�Q���X�7}h�5+���9�c���k;+��"�$�7y�č�-�&��5R}����\ΰ��2tW<#�c��@��U,�K٣��4��i�`g2{�@,	���I`�
��K���#�.�"�%`�R{\���q�l�.�_�U�܅$���Xէ�P N�gR�����:
�������^��QN�ѹ��Z��}���HMR���=�,A:5���m1cp(F���}5V�{�:���a|��JeDh򒣛�Xs~N���̔M>�����@$�p}����[�������^�*�Z1�R�3���7�@:�t�E[������X=�0�w�T!9��5�ܬj5�9���D�u@���@�N��j�1..v�c��]@�A?��v����Fn�UWi_�S��ۜ�w�zw���[�Q!��e�gP-����霃�4�dKmJ�v؊�ޥhKW�?j�+�&7�i5�� �s�I�o��d�o�$*�Ã��j2C~��0���2!�T��YZI��EG�J~�fAw��r�[�:�0U���Vƻ���f���ʁ.��t+:�d����7�*�'���&׍*��L� �T�k�әщ��P�������0J�'�0Yj��@�}A"^_��"�}2Flu/վ��r4L�kz�^ނ���Ϸb� �g[����R����M��^�t�E�R��Tm��sӑ�9I�[� �u�%�9)w�i�"\�Õ
w��j�D-4iht�p�S|���7ܳ_�f���=�̀�tt`�=�!�� qU����[�D���d��t�(2�r�F����S(�z�}���ȴtI��l���h�Lv 2��C�@��e����(��_FPU���V0G,��2y5�ؾ|Wz|��p�B�`\����������Cm��	N�R�':|�U���J�Լ�@߶wz��WQ��ehÂ��U&"%�n�i�D����R�50e�Vvh�?�ڢ蛗�k\.Н
f
�(Ρu�_`��H�~K�.Q�6�C�T:�l$�*����5
��.3~]/`�&�v�G����� 0l
��m�e��g�	�����:1��,�Orw�_O(�!׏����b=3���%�_r-zp��GS� C����s�r��Aj7�"n��Hߣ<ȳ��n�d�
P���n"��4 ,8���4��C�?��A+Mbk��CU�aɲ�,��"�ʊƜ@�/*귉)�̆�_Ǻ;_��6!o,���t��`#z���쉋I0��0=o����;d��W�W	x�B�"c�F=���AH���w2�{��o�u����(�c�B^����l���ʡS����0.D4ZC�~���z��K`���2
��Za%[&���F�I�-w�gWy�c'����7��`<�uN�	C��D�o=_L�>D��"�YZ�?CG�O�/5��a��7�1'�g$�R���5y�q}쪜j^R�9V�F�X���x`4��B���g�1EJd���9^X`yl��U?R1Z�o�n;3�ӆ4��E��L��� H�(Y��U�6��_�e��M9�_0Y��cx!Wq���I<�߸��y��]}��&���{G�F�w�;Vף�<��|��6�ԩ�-[S@d�jmS�:�Kdt{��3Ӿ��f�K���oOi��$��P%��~ �ju�$�̌��G�C�nSoS](�`����ų�j���1R��`>�2G����Ö&�H%��U��(�|!L��;�����j� ua$�n�΢<'��t���Y��c��������Y��Y�1{F;��.���:��}��9{6�`�K7� bJ,�.��+�@*��ج��������V'73}\���wN�z�8��_��9T�}���Z4\VY�������be���Yn	�e�z��}D��������ǈ Ebi���1-�/�@�
�g���`����M_S����1�r�/��ы�:�d�!u�?&�Tf�sM��N�Em��k'�3e��ͻ�c�N�2�ٴ�Ѩ�w���3�i'�.���a�����Tl-_��
�ٙ}��u��bX D�9d)����J0xm���H������+DZ�c�*���|�Tm�ڀDCT_�J.�W�ls
L��GJQ8�^�p�{��ۆU�W�@$Kne�4��AMJ���$�|��PƼ���z�S��I&7�ك�@�!�q���2f��[���$˄Y8*
o�*?���&�)��M+[�&���E��.s�
/���zSd�W 	��f] ���:^I�%�m��j��r����Fi��$ w
�V���m4B� y��0|��J��c)�5Oe���Hu.�ۼ�_�I�yr=k�mb7 ?��@>�Cw�j�O�<�]Uª`�Ԃr%�1W~K��� c�`O��!�����\K&z�o��K�C��])�v�ru�Ϸ���Y�&�N#@�+PSÁ��e)Pp7�v������P�'��?_ߨUW��OJR��.�U"&��1���5�B�*�U����6S+��2VJ�2N��C�|��(7D^/����s�3^���㵁}�-�X���(���!]�׳�����&���	q���~|8)Eƥ@��Ua��8�:zr�4�m�n���B(����Ywq�$l�j�q*�o^��K1�!g{7~1�̛�o�L�����#�ĸ�F��F��9z.Qɫ�p���!�V�	�f��U
$_FQ
p���Nk,`k�a�L���>^�A	nVろRF���A��i��f�T՛�QCj
���ĩ�{�ʉ�C_�#����7{s�����ǪCe�@4�(��l%M$�VCS�O7��� � Ŀ|����"�Kl�)�I4�~�"�G���U��v��$g�l�jr3ev��Ot��v��(�-L�Hv�����<�@�SË^ѽ�ro�B7��n�g6,UK�In��+�t`P����"A�r5m5)��Z�*�I��	�-��ha�â�c%���l#��v�}Y03k
�+�Z[���^{$I ��;/����w���A��99�)�S��l)���b�m��Q��3�BD�2�~���F��P�ŘbA�D�3>��)G���O����"{��a���W�Ĉ��'7~ug���/��O�]^š^�8����0S£���D��{I��G����LE��Ֆ����@�?U�+�b����rEgj̈́������Ȗ��ã�Pd�W��z8�p2�G��*���sg||���y��ֳ��%�o�#7Ů��,5�gp2ϖ��,������SA��b�;S�r�V���o��㙗R��+&������]��ɱVו����e���B�:��@�I)����e�3�Q��|�B���NY"W���sŃ��r���D�ـ�ɬ?��l�g̸igl��O^z�^"���Y�|8Ż:�����*�`Y��f�i+��<K�=4�<�
���������0�@[2}�[r�j�#�5�D�MF<< 6�S6lM$-�HC�N�$φiJwp��h�7$\�,��x��]^t̖��"/w���<n�>�u_j=߅����Ā��wSpLQ
����*Eh;�,D@�� ֦�q�Ļ�ҋF>�~g.w�?�6v�����I� �m%0w��[����[$[V5�5Ba�>v�[�h�ї*GŠ��'z�˂�X�^"��e�^�uMߎ\3�9���Bp��嚟�7D �J�Gxw,�v��l�p�l��K�C� ��: �I��0o�h^�	����^���_��ɵ�!��@�Bs.)��	����?�]��AP��H� ��f�����9Ц� ����1��(�A��=���v��ꠄ���n%�t�pZ�?��&A��E6�+�b�$�C�}#Y��!�咤<Ų�)�s`6�SD��*�D+�ZV0�u�B�OY$��45����y��Y>�_��<J�), �O��f��Dޙi1�@Yς�=�͕�|/�*ujN�mF����V�C/�VB���#�fKU������n�G����a�	���r7����Y-�9	�.-�͝"%��
n�/��W�puMu��::��>I3I2b�it�^��ps���bfp�mE�ϯ�0v��D��� 2�wmW"OT��	]蟢kTr_�	q����z����^+5ףT-~v�&�x��TXy�'�u⠱���=,^�`g�.+r�t��q�m�pK�c�[na�񓚪8�[o'q�v(GR�n3���U���pG����*����ѱg��	HP�+��b+vk!��ߍ��Cj�ӓ6�Dћ,�E��	#�z��Zbd�';��#���spJP�؎�R���D(dj�\��+iM!��&��-N7�+�l��o�c��{l�-W�� �{M:8E?�N�u�|��G����1��g�D��0ƭ����i�ȥ\�ǹM܃hu�Q��N�ġV��4M���!O�i8�l�R���&@�m����(w���JU׶���H K��$��m�B?��[�ٔw��#J�-G0s*E�����G�i� ���2j~FB[��T��(+�%H���Դq����23ar�c>2�z�I�ԊN����.�د�]2F�l�`ЅPVB���T��ƺ��m�L���e�q��.��T��n�]N�b+DZ����'���U	�h�Z�w���ٓa$�ś�3Y�Ő�5�������P�קt����릖��\�kS=���i�ުdC5�zS�F�����l���c$P��Ӌ�%#}���$A�C�Ͽ���_�ۘ�!�����%`����Ag/�@-�:A�p��ȅ�V'�x��7���o2iD_��I��?��;��T]�H@E+ZK��O����m�9Gdܰ(�AȋK"Bh�y[���׷l3��M����F�P"��a�v.�\� �ְǩ�G=*�q�H�䲀o�E��.</��B�AÞ�&C�1�i�`~�������ꇺ�rQ�g�.�!�\a�l���⾃_�K�JD ����$�#�M�������|�+�Cd���V>*�������\�F���p��~>��e�|���K:����x@�QTzb�Ia�{���s����\���ǉ�������Gi5�+y<2L�0!�a��B��X4xC|�
pJ?�v��xV#a�J��:�G*�|� .����L_�cW��ˁzR<�u7�u��vS(�V�y�����U�O��T[6�*��eJB�1������X���bȁ��H�-�*��'�˧����T�4�l�H�<D��p?�2�B;�~��#��cǟ��)/P�=�ʈ�H�d𛭃�4Vz_�ma_
sk(�S�Ű؝�8�M��~���6�AH�MII�Nȡ�6����M)���\������w��,h0	����0��o��G=<hT�Ml=�PQU/C*��g>"�r ��M���a^�T�����a5V
��J�DM;B/M�h���W�8�e#��6G�P�A|�"���<�셥^&��!VS�fג�A�?K�uv�Н��~�E6�?#��n!�`�+�����W��Fm��b�(#Z���[1o��0A�M���96"��Z�7G6�b*�qG���ї؋Wtm�����a�%�n�W����#E��mR� �`8ssw%a^7ǵY�/��N�Y$-�H�{��I��[�-�0!AcPtr63�(�����s&���7nH��^74u ����@�Y�P'f�����:}�m�A�� i���G�Eҋ>$�pC��eic���Xq��kE@�l��L�x}�T���E~��9*��CD�zyyg�b���u�5���(=�vS��(a$�O�}�wp9��M�T������ �+���\��	K�1U�=Ȁ[�F�o>�M(�0o�m���V��
>�X[������H���1d�aٿ1�{��lP�ҋ�z���ox�ۏ̆cP���G�5��,��gri�o���u,aѡhs��nG�&/�Ĉ؄��>�X��`?��)�=�dfqE�|c�#��D�-Ҭc�0X�/]@�2喘6+�G�_V���>P�@�uV\�r)Q��!����п�`���i��Y^~��W��<iX�Od>6$��ҳo����l<B� �~����������6���XU����Y�.�i�i��ja�FKf�A��@>�V����{��th�y.AV��k4rh2O�8̾�oq�
�aiMfun���/�ijͣ\��q���m��b)�5G���ɚUTc��3W���۾z�Rn��~Qs�̈�����l�����B��F�T�n��v�-�n�L���d v�@�9&`��wC�8��`q�$M!˘v����MF�hb�Κ5pѴ�p�Ԛ���?4p-WquHT�y����~Q;s�V�KW���׊�c��c�Żz7�Z��������2"i��2�We@��Q���F/X�(�	U3J��c ��vң�����G��5��K���W�o�5���?J�T�k���Ű8nd�i� 
}T���[�t.~߫�F$��pϪZ#E�`�b�ŷ�)Zw���T��̀�Q��~�@�xw�O�B�&.�"��+��`��d�B���?캻B*	!�Q�}9�[��xԢ�NʉG�߳3�}Ł}Sd^a��.q���:�Bov
n���?�+G�ƴϝ���:/�����+"^	p��lN�?����mW�N�oA�>��r�ЎG`Ʋ�Z�@�.ߦ�J���E�������T֢��:#r �[;�Y��ӷ� �d �7�-��fղ�J�P�v��PW)��!-0�m:ee�ss��7���d�����X,R�u�P�C�X�;~������T��y�j҂N��%pĤP�ZD��;�H-	����e�b�����b��h�*C�Vh��Z����_y��?���\��,v����Q��:�K3�񏩓�*����"��1�}E��iӷ��/��wu2*�����6���C��X3a�YO��MuO�-R�Z⬗#�7m��
�q���d��6#����y����z}��/S`pK�>s��%/��D����$�-1�cQ��r3A�F�g�8�*�l���)G�,U=��������?�z�f���ɱg�����tꘊ�[w�g�<�Ii����$݇u��S�>𠗥d�G�͖�W$^�V���<�*k�4��@��ZR�t�u[�0{L+��!r0~<��J,�_����بz�'��K[.td�oe��h�L..����꿘S��,@~����N{W8%B�::� mj��?i9U�0G�ωG�X��Ia73&��t�D��*ަ7?��2֏�[��]��1b�*&��@;��:����IcB����c��A�K��߰}�睚�����q�����D����8W�{�Gg\~;:���9�<�h��W�,�����Ye����;IV�=~c+
��+-l��ʜC`c�P�b͘���}T:��cRQ�?���sJ�*́9���D`�0�N��fm����
S ���^�O�9Q�kT�f�q��m�cu]zq�2�*娀V�.������*Rr�J���J�)름>x�/HX�m �m(⟡7��s5HLr��$�u��MS��̀���{"6q
ϰ�m�Y�Wf}�5ڭ�������+@^�p�KM��*7��Ɠ����܋v	��) y���7��b�=!����Xx�����M���z3k��	$��	/����2O��!�I~��I2ٽ����*;ǋ#x�g5Q䒞$�����:j�{��`��k�)qh�{��o������壒e�����?�c����W�)��x��/	�'�QZ|�;����Nf�il�� lċ.M������Ci/��'{�9�>{��`��Y~�E4���[�����U`?�g�X+L8�6eP�_L�yz��'dZ�D峅s��B╢���$K'��BAx����F��o[%/�!W�f���݃�[�}j��I6V�yz��E2:
Vj<ĥ���O���cX��:���)h��H2�
A�h��6���q���p��M͎@]�)�D����1z۴NT���P&u������7r����!����D���q���E��Gm��܏�YTEF%�q���o'��x�($�^8���a���m���}��<�,W�{�Jp$̚� �W���(�D��fsn�%o������!���1聱-� >��{�M�x�3N��L���˳]!��RɨV;@n�E"����{k�V�7��ܚ�4=���GgJ1���˜�4����v�f��E:�=�̱=q��z��>� dv���`+�
�!��*�}��$� d�S���=��Ҽ�q�5�k6��,���@.I?�T��
�����*ҧ��� dtaB��5�aoB�Kpa��1'Kbp7Kj.��gg�T�_�����M5��?H�K�����RL��W���
�M��P�v���h��$��\m���ӓ �`���ǣ��ϐ�ɵ�k��G��"_~<�����n��Z�WIG4�q?�d�`�I�$�r&��Yſ�6x���x��P��U�a�e�Vo�Y/(c������V2� �������.]�p�9�ͺ���Y��S��,�k]Im�.ꕖ�ɕ�s`��"�T�M0ĭ������]��(��=���j�&с"�j��}PK��{(ͮd7�U]��5�%(��`¨�
��k���/6�*oi����;�l�.tO���L�602�r���ֿ�|����ec��!�3L��m�`b{�����������xIG��ڴX^�Z��g6H.��T�f��!
'\��LO�M&�1X��}U��7��4Ya�i��Fe J�߸j���6.�l=�����C�U} ���^�5����;-b�3C��@�5Iް�?]/�:���*'���l��uVL��{YXĬ��}��F���k[gp$gq��E�ӯ��=^�G�J���6����w&�f����8L��c�UJ�ޢ!�0>�57?��a[$��+�"E!�ҽ�� "�v��Δ��V������t��@u���:�W�٫�Ш"�)/�q�	�ՙn��N��p�2�S�'H0-�W�ި����^}�t���f��h��wb��0f�v��Y�X��F��j`�_�2�3��f� L�
�K�A�Y���y�c�!�eL�������3H؊3a.�ćpt�N�ް��#�芅%�i�+���B` �&,p���@��	��N~,�U�kS�i����<��M���Qx�Z�YV��}����}�򗝱�n��`,\�e0_ܹR��y8GB_p3��0ƅ5�:�ln������͘����O5��a�g��`Fv��W��GsLs�`(��42�$���o���Z�rET�-7�D�8�G��t�J?�H1f�(K�>\����v1��8�^��u��6}��a��IDܤQoxJ�N�y�:��˚a�X� X�4R9�~�P�����O�#>>v�[�c��)�t?�/O�8��b��U�o`��dv;����
�VI 1���d#۱�|Z%�9r�o����i�u徻��·���-J�os_�E��EFg34/���ٱ2�_I���ր���ߩ4������;9��T��Y�ѯ:��<pw:Rz�=g�\�*��a�����<K?�๥�3�⧛R�;�R�*_�@LDc��>3,xh�E �_����|�Gef{eCYqa���&���6����y��w߂W�N�H�n��ݎ�9 �� 0AX�ǁ9T�L�봘���m�@y�0J���*f&s�-QY�/����S^-��<��j�+ȒLѡ<,�1:%m�lJ	& �C����h�I�zU4S�~�%_+��q:�ۺ�8�XЇ�~���럸S�x0�Gv'0�i,<�_��H�	W�����%��v��@�'�Q�\>u;_�swF����gF�
fo��r�xeR���Sl9%l�ݮ7C�3l�a��Z��?��c~_LB}"r�N�U�P=q��]���H�t,]���L�cJ��9{�r�Y:O.X mO;9"M<>��{:o�y-�^* ��#s�*�$&t��.�*L���i��Xw�,o�a�M�6+/keg��p׮�7���Rc�j�..���׵���(��N� �[�� in:G��I�q5C�N<��=Ә[������P�hz�m͡IP�b��@Î�ܔ[���4!�g0R��o%�hk��Eݚ8�WPe��Pf�U��@ �9x�UOIsT�OW����f��B�C�Pۤ|앣��y��!p�Ud�g��2liDG�����~��C<Z��S�������xO��;���A����y9L�Y�S�)�B�-;ɐ�55E\�X�j{i?> �b��+A �4��H�f�uk�O9g��߉.�w�
<֩��Fx`E?��ʑ�"X�j1���Q�:��a�\�>���<�<Oq�+
޴gx�C�a��|Z�`r�(����r�	z��?�oxa��3�ogy$*r\�>E�厷�]8��\���ƚ���Dae�ƴ#6#\Z��g��/����)�X%� �9�5�����o�T��2v���ԋ�`�F�yw����:8TG���/ci�$N ~�{�^�ƿ�}ʝ&R{D1�h�� 5�.bi<�hb�5%�Ec <2���u��B�Y&�����@z$j>�r���{~��{����kZ�S���}Yc���Z�#��E��w�e6�*qha��S�������<����4��>�fK�Um7c�[f�v�3�#S4�CA�FΪ�/~�:�AW/����W����j��c�A��0q�ĭ���_�_l�a=H��IZ��/�n����9r�F6/��o٥���UoTR-3p�Ԇa,�8�qzO�����	=��'�%|ulB_>у�P32u;�s\��.��R� DE�ǻi��w��b�Fa��<���홒��o�3D��s@� ����PI��s�bä�A��I�~Wm^�859+Sg�����\(U4���� i����qNk�|������3���S틛$'#�PE�w46$7̃�|>�bˆ�!<洔�p M!?�t�F���V �'ە�#XR�%�n�)��z�_����h.�i���a��Y�K��9K�d*��N��������֒~S#R5R�hk!��f|/q��D��v�h�[p��}�m�=���j�$�v8�%u����7���=���v �:���]vܗ�����`E>�`��L�m�����'�(CD�[�$���3�3�o�y������h�tr/[ؑ@SYw�k�^��}�\<����d���>��m�a��X��W6#��D�n��g6s$e��,҅2���aD��>Cq� ��gB����y����`�N�r��k� M�D������$�5������)��c\)�������mA�Gar9�>���v�}�)�h㒂f�\ث'U��l�B�M;�Z#��32o{��.u��;�3v�S�G�)p_���8��G�U	��h�*���Y\�wtL����鳸�J�,-��ڧ�8Aht�8�)�flzcH[E7끸=��R�_�X���~|��JY�=J�3(�E1���핟&�w��gi_a���'ʓ����+ވ����]m{���#�b�X��\%�̬P��*C
nC.�e4�_�����7%tmsT��4Z�	����T�f�O[��@,La��&?W�yd�RH{�L���(p�d�r���?�}�e��E/����i�E�# bY�M��]ՙ�}%ܢr��1��-�=�<Կ(�N&c�e&RC}�sjt�W����C�Ҳ]52{�$p,����O�խq��܄H��5EY>5���S��ͻ�%��\�,�뽻�?G��1Vz��%@�j��>;&��R'IN`,��f[�#Pa�Q�n�(�Y�ҿ2�B7�i�'���	�'��xz�_+�Th�B�@X�U�.��*��:�b�M`������	#)���Σɹ���:��k�u��&����z3d�t������!Vf���x���o/�ۀ� QL0}���Ŏg�zt��1����@_��P��X����5�*��|�� �w�?PHA��}i��<e4A��m~Ѝ�J۾3D�Ը��G��ARͿ.+�H�U|�ak
��;m��O�3`�5S�*��@�HR��D`§V����'����5��Q�sb3oJ�e�Q�d��D�Y���h�0J��AO�6]0�����\���:+&s J���KY�cEI�/,ƴ�}���#IUd���_��Ū�qg�g�	�\��ю����� :^X�������N�
Ch�=:ҵ��
�)�-��'�q2�S�C)>�7�4.���5�2���s��/��Fk��U�6���Z�C���*��+e��n��`p`[l5Z"RҢ��"[�m�oK��jruP�Dj��NU��MO�~�$&�]%�:gWT"1�9�*��)\-�m�&�8��!$��ʢ��GiL#0�%y�>y��E ���]�����v ���NQ�q��$��3��2z�w[��=����jm�q-az����!����j���<�R+�'��j=i@���)}pI##�c�{�â��6�c�x<�9���57�Y5�	��Ѥy�ΧRh�[�:�(��c>��m7��]>&���n�cҎW�h=_�mti\�a�c>����Ip�:%i�C��rP�!&�֮��䖳�33���"��@�?��5��1.��A�?B~�rD��3Ou>�Ulr �:�L��TBo�l��b�����=@��vՀ� ��!(�.vjK�����l�y�sQ�H�UvJ�w:KG�]��+-\d>�VoK�@�u=N�F-+Y,3$2�H��6` ��}��o�ɽB��%�@�2�r�&x���̆`�|�B_�B�.��S���=�F��c\�v����?����K�tc>}ݜ�>�~Zz���}Mp8b�9���ꙸ�w{+-���z����t)���{���d-�j7�zmw�Y�����.2�~��uD���]b������,Ø�cG�hQy�=�+pf���E���Q�2�4�&>o��"�$�6�K����B�ћ%�����Ķ�p�����o�Ez�@5�"|L�:P��zG~5�M��-����}��G��OYe� �@B�X'�����j��`����(v����4�NP�J����Nskݬ����h�vcޏa�ʯ�~��SJ��yӥѥO����#����@��s�3Oɥ/�M��N�PHUL�F�I�٧�1d/&�W����eE���T�
{��!��Jrbt��<2ܨ�{�����)�DЛm�/�aц�*�����ҭ"L
E7��7=leKV����8��'�p��/�kNK���bI��FM��$��o= �
k��`�a:�������������e�
j2��������韑}��,����UZE�0���*�Y[]}�+( 4Ь��lW���Q����?pp� z/�$�����8o.N��𫐯� �Ɯb�l�;�n5\�D;��^��o�� j� �z�7ϟ$�C;�T
�ȅ#'���P��P�S��^���<��!]�F%c�O�s ��M>�*��� �$?�9U��菺o&��*�D\:4����P
�7&��X^���[#�S0t䷑�|� $I��C:�f��\�^I�/A�pA�n
$��gyL��x�ߪ0��'[���}����n��g�'>�* ��.R�����x�h�Ö�_0��Yc�>�0�E8G��8~ ��i3{RYe��Y��
�v�s�赬���Am�#�ͻ��N�+�u��s�鰗%
�<|#�R@6�;�Dief��!= ��l��� ٺ:I� �n�q�R0�i'�w����?'��맹�,�2vZ��P�|q���Le@���
i������M-�Df���P'�Y�У��:���lG� ��/��_ ����ŕ㫻lu+B�6�9GEP�&�2����+í�u�1��/�q\��7;��	���Ի9�M�ifF`�}�jŎ{R�� ����,�Ld�
��\#�ݍ�L��#�HcSǭ۶���8���M��4�}\��lY`�6<
y� ����nF9Ppb��ka�j|��ra�������<�p�ҷa��R�͗��"4��il̈�0����V�˹ uN����Jp����f�ߓ�.}��৲�f$u�	1���Hd�����G/Q�k�Ͷ)�r��b�Ę�I�b�ˣ
m7��S���J����de�㽟�>N���C[N�"�\�B ��'���B(�*�N� �L��nH��$l���I;h]��Q������u�E�y��[�������JI\J��K(�����exm�@!�d��N��QՊ
_J����$��
A��L��Ѧ]���5���*���������u��@��p9�1,$�#�KDPX��W�Թ��k�ݏ#��.�������̝2y7N ��]���������(el"a�����G�I���[n�*�J^�_&�����?:Z��:��%�1�k�3��(�&'�f�z������Uds�wt��@yڠ6�	�zL���XX�qT�W��n$�?�TԚ���!�F/�ء������)��׬.v��w(��Wh��9���\���a6���$�S�� ��H���Ie���g��C4�(��<aZs��̠��#�K5�+;��g6"L9�iI�"+`@,�0��8��"���	Xm�Ьݔ�� f�o��Hd��/=�J�<1�;V���Z���D�ؓD����ٷ�������=�a����%bA�,R] �N�E��r��l��<!�m��ID��!X�&� ��ךI�*.\�.�b=�hv�[!,Lm��ʳ�P��� ��1v}(�Y�y�?!�I���+Ѥ��z�=���X�,�'z U)^/b�+��zǙ�m;(����8�d�53ىz{���� ���bV��^�3]����LZ��L��H�,.�����nITD�S�^�G�R=�Dl�Β8�Z����rR�"���i���R�+�ݽM3�^�Q����R�w��<R>����)d�_`e.k�-aS���Һ�> BWH-_���0>2L�Rr�l��X�-�������S��� ~���G��!3=�����m*|����r,=��.	<n�`瓵Զ)%��U"�d����	@��toܨ�>�̈��5a�V	9��}1I��K�$�Bw��*h��6}��o�q����r�c��S(꛽��V+��J�h�]��z�Bp�E�a5���ߤ�r4�ZN5�� (���7�C��t�*��:�x9����td�|]nO�M��`�ҥDY�l֯����߽�Ď�9�?�Y�U�FV77<v�x�M�(.Ʌ��v�-�������Nୖ�b#ew�z��(k.a�~��=���9�>��2K	�s!l����-�䜮o�ߌ
�� � ]`�M*�_���qv��"Y^ubx��f���$ϝOAls�T����>�G(Ӡ��+��b4���K�od<��_?k�փͼ`�Γ�!K?�����SeyhdsWɺ������r@�r��e��ZՔK��
��x�@�� ��%AP+�YR\�� ��ȩiv
�ށ�#���?���Z��V��lr��h/���[�uV�`h"r���8"a�A=_��)��K�e�?�lio}.�0ZUك9YIƧ�맮��.�-��&;0�ZR�dZ��T��=@(H`K���1�,�]n4��Q{�2�g��]G�҉¯�#�����L�?�|�-B�e��2�^�`�W�n��	���O�#)��/����v��� ���hcx_��`F>I<^��	~�֍ʉ���J���[��]����f�?��e�'a4Q��@!��f��-����b'�؎�WBn�K�ش��̎���
���(��I���
*͢������=�)E.�Ͳw������!�

�4��8J�l�����}Gp7�P�d���{汲O�7H6���_(�R�hJ�j`J9G�e��d�;K!N�K��.H{,��׳ъ������ս��g�7e��q��ܱ�"�V��\�C����}�`�n��hŽ��αҟ␈����4N�B���c���)��?=1���%�1������� �)w�=�_K�s�x���WF�S}_��/�	�����`��/M�0֋����W��0]�H�nr�l�Wϻ�7u��2<�7����i#���xˤ� +���(Z;�3�� �9a���*�w�Z�����:��N��!ߋ���=��w��`�`��'憊7�C��!W)��*?J�ߟ�fK
Ҫ��7��,����n-$�-�PC7�� ���7���4�ͩ���� ]3��Gl���s�����(^m'��5�y�Q���tڄ�G��� Y�ǯ"��v@�Y�$Pl$�zg�Q��/-�����a��!ʶT�'�4�d��[j�ᛉ��{c�H���$�ޒ01<;-/���e�����B��ptY������&sU�w��:�'^��D=X���p���V��NX� �u�+y~�HH"̍h��pF\>�]#��C�P�F
����ؒe�\�����JQ�5a��W�Y,hIA��y������J�z��g5�˰���^d%̲��Y����j�c���"C�7LY��;k� �|�tH��"�c%�=`��R�em�&����q�{�B�C���晍W�39c�Z 3V�'Ə���f�cp�rb�vǬ$�=	��@����c���a�ΕOkt_��`\�g�ZK�u����%�o�l�)Eu�J=�̟(J�U�\�A��<
�CTJ�u�����\�Y�=�8���{�g���d�(�+^����j ���ӑ�9~5H0���Qu�f����?�N�%uA� �>߇Tέz>��D�3%;��ۥ#���_A���H��y����#hY��]:��J����|��|øp�"QK�b��1���T�qW0@��z�=ƞP�%_"��F� ���Tao��������z�CEns#��E��$����¼���!G�d"C�w���]��6!�gٕv����~ڲ�Q�y���������&U1Xyl���=�a�j�^@���n���%Ƨ]n�5Hq,|������h�}���S�l�*�r'��^�^8��*́��8(K��d��y����Vϻ&"�M�7`�P�}i����CT3:�Vҫ�W�Z8bB��ݟ��ͥ|����-`�NU�!�R�1E.i֜�������#������c`��)*��$���R��죐ol��m-���#8�����N������� ���vlFP�f�wz,`"Q�%�z�+���Ya�1��"�'�^�OT]�����`�Z����m�B;�	�P�~�/��ŝ
U���(A�5��λ�X��/�;��V*`�a!�M���e�O5dF��c�_c�D �]�����_SVw}���"��	�'YR��z"�J�"���{�������;R2�)&{�JK�/tH���\7=��
�˿��dad&
�#!:�,/�;<ώ� f�p1UC�O'�=#n�/L�_ԝ��x@�K3Z+]�R?���@���SO��~T�i/>4�L�|�{ْ4�����kN�>(�Z6�$�[�S�l��/x�'���H���N�k�kÍ���ANO"��\���Ŧ[Ґ@��E���O�t4֫�<.��5����J�Ӥn�E�^���}��ri<����TYj�Սz���[T���dZ�����H�]Ƣ���w�'.����>6�c��m(�s)���[Ͼ�l���̤Z"��y��\*���!k�0y!�gUm��.��H�IQ����`��]lz���?[B�3�J���q�~3M�����4>7T�b=Dd��"ȃῙ�v�'Y�0�6�����4ĨC�.�Ae��<���UMP1��V}ܾ���YM�c�Z9	!ɰ�!Ac�خ��m[<CNt�&t���b��.|�� "��:��{lo�7	����h�p�k8��H�CƔNO����e�#��{R�<�����h@)��^li&�Hruˢ��ޜ2����nb���;NI7�4b㼺X�ʍ�K	�/���V�7�}΀����Uٴe�r��:F��
9��ſ`Tʅ_ ��GΖp����h��4L�]�� �kR\�����SL�l!A��p.gAR
r�K��a:g���'-�����PKx܏'�7��Yt䜶�&q%�!>Td.A����{r�쯽0�](wJ]���^�m[�;�uJS��n�}q�a;�
���~������}��V��aP}8�	�%E�J�[��b���F׶�d,����JF��<�}�K��Xo^SB���C/�� WJ��$��{���o�izgLp�º��JƧ�>b�nlo4�*��V�^�fRA��G����-��D��i��v�VW�(�(�! �n��º�;���Ȫ�v���d=��W�,��]�o�DfL��,夋3{�Ib@����\Y��׫#�ƞS2��E`BS� K�-U蜁�k��1`�124����*���-/A�>Anv��󔰑�s���10�m�>� hA��A����:���țaB�Og�Ud9�mʸ�-e�ƻ|VX*JD� �D�z?����3'<k�3�['���	,+�И����3�GD��r7�q��F{�13$&��Ji�/�^�����6���ոD���5
F^yX`��2��_���p����?a����0�s�MۈrĄV@}����~���4ڙÍ�A���jlm�� �Z�?��!�4pD�����-v��m,ё�͐<��͡\sDݸ�<��A�%�9��������i9�Lu��;��� 5l/��hh�i|*O���*�����^è�����;5<s�F��ѥ�n���������X���.������x�+	M����uO�1�d=ڂ��W|Ou��=�2k�0�H�C�ܰE3�rr� ��\�y\%�e�%�6�s� y�xL!l�M2D�z
��2��d0G���jh��[�P^�/�Tw����\�r>���#�jf�jk"�����PUO�1UC���T�|�K�P�����W2���Q�X�(G)Cg��.}iyOd�:�6P "w��V�7����_���֛��A��_�r����S(�<� UE�b��]���|��(�ٷ�@u�҅-? ��Y�`��Byh�Ɓ����"۵U � �m
:�yb��� "�}�o�|88ڀ�d$D�W�W��d1��dU�����$g�Ôɤ;uv��bu6�H�X��=Q���~!.U���Z0^$Z@�X,|+����_k���p�������;)�9�vc����lL�ݱ`s^BD��ů�)�"�h�����7���L��bY��v�SHc6k�0է(=�LĒ)��x�*ܒ��mkNr�8��?��� '��y�Vqi�J�ʻ�u#W���A���wƹt��������ПeC8T�dO��]�#��Ȥ$�ꬼ�M>׮�g�*8�$;����A�����įl��XKf���^��?�cZ7���*�)����/��թJ���P�Ň�U/�!RD���8#�h~��N����n���W�zb,�2-t�m�A�.��M���7��ց�fŒ�x7��wD.X�PiTuh�v�(j�53��?G�=�����������t�F�>�y
�8�#�$���K���r6&H�g�����?CZ##��n����a�y�T� 9	��v�;V��?��2P7|���_���U���F���H�E�����l�}D����I�� L"8s���/��s���z�)��n����N�Se��D�w���L��؜].��K��;��{��'}�K�?L �|1 ���I�W37 '�:G�g?U���$�VPl�Pb3��SX+>�0:(��O8�X��W��0= �	��g���m�9X�@.�<i���$�z��A<��r-��%M@;��nE!P,��e] �b����#�"���,��\�k��I�e�.#|���TD'�~�8�&$�n˙�:��(w�=���� }iuA���Mw��k��vX�;bg��d-��256Ȓ��c�����#��ױU �.�}i쭋ֵ	�~�63;˃��\��S������a�BfX۬��~�.�P�
��z�����q��h�SY��v�c�!��1�8B�|�>�z�n�%�B �:�M�Mr��v�Px��f�a�-c��w9�MiF eb(�6c��f�`-%S@Fq�w<�4���n���n�ʰ{!��A�7��fųi%42%�7=�u�d�,~���`T�I�!�H������LK5������O����c/t��c0��V�b}�^���N�	�(L؉0������[��gYH����jsĚn�T� q�Ңd�o0�N$(�F�a�u^��7"���
��k'o��1&[Z���uȽ��;���� �Gc�Z�e�>�v��_��	�X�����'�,!iru�Rr}4g��8�op=�:Ӱ%�X�h���0�M7����a7�p �>"%�'Yg�w.���" !{2QT�A]5!�|7Wϐ~.�@Yo�vR�^�#�o�*SV1�����ak`@�c��:�u��p$�hB������&�T)�U�ٗ���;\��ז��B��&��@��y+"+�~�^l`Z���C��݀"�5i��t^T`k���/�� =��?�͆N8H,������Pk�fm�y a@���᭘J��]�2�E�Mgwf���|�t��,�)b�F>��M,�-'@�<	& ���a�n�¥W	�����-����lg&Vn�z���}��r+e7��#�{�w��R�`}
�}�T��y:�����Q�����P,��(��績)N����S�ύ��l�kDOi��6p���h��L�U��W�k3�?�PX�m"����B��giWoϢ�wxCm�
���j�-z�?�HUQ<T`	���b6B�M��/Iޓ���jۻ\ݳ8�?u�\�k��C�1�ay�d�3pּ�;�R]�`�%�E�1x!R���s�r���X�������E l���]�h�N#�l�B������a��N�r�&)�[$��Y�.� Z�������t�Z�#L�u>��X�%��M���?�s�p+�>ΐi�m�(yntK]�+h���Fd{[��(����D=��8w����̓~p�4UB&M��y��B<�_�~,jB�KZ$\l2�.Ld $J�*�$��f��.ñ�/���Y�a�t���A�,�W"�����<�iK�@煜��{���(���Y�{�B5����N ,��V�H\�4	+iY�������Ѫ{GlC�N��'�.�����R[������S�-���؊�V��+�u|U��4�d����l�GC3���RP���)r���~v�9|f�~�b&n�nV_(�[�Vyh�}�6z6�~��:�rr��CF��E����;�KQ7U��-ag�\�䎞�d��$�� 61&UWJg#�\W���z�C��Y�3�����2��sZ����fO�zو��Q`i؈��MI`*O��<�s�?)��A=��U�&�����|i�Z�y8��	� �z��AK䧞�,�A��2tHT?j�bc�h��(d��\���Ë�i��&���{P�Xk�(�>��ZS�����X�`��ƪ9� )�+%�Vη�=ʂ,���7}�Y-�O^��Փ�z"��ez���9���d�VO���R��&�"�!���"�Nd����
�M�|.J���E�F�)�>�4�L1m(�����U�a��d�SJ?p$�R:�_
 ~�����Q���� ��lb�8��(�|���V9���4��1a�rV��ᵦU�[�@+��t���O����rp]���y��<��#
���T���~�z�9puI�W�Ax�p�_/����(������H��ρ=�j���l"Z��5ɰT״v��9���-��/����Y�ɯ]˦�C~� E-�7�ȧ�/�\��
/����8N���1�:{D�0��
�U�[�J�򰵦d�C�z|R`�*�&X���#�83����$�.�y�e�eɌ�)N�sS�n�|5�N�����1�-3Ǎ��Q-�J#&�+����`��p��W^/l�Zg+��X������ Y*~m���}h�V���4������W���J�F��u��6�5~�HՆWH%�4;{B@!�;^"�~�$�=8��vD!��=��ɭ��?���ךUr��5h�%W۩@���>�R��w8@���C�G娱BI�|r��[��d�{-�*�mo]�V�-8���L�y�Ǵ^_YE�F�3�M�M�i�t�Z2ط��h��`,ۘ�{��J�@�s��,��Ȥ}K;g\�!���aў���u�q?�>�u?y��k�Y�1<�Sx .�������ǘ�T'$�H���CɁ|��!JG��\�'�/�����W��n�5 ~H�ú��lL���P@n��v����apq�ϔin��F�J��!���$"Ƿb�t��<�?㹋m�:%ă�l}KК�;��ۍ���{�nD�m�|�7p����)��K�4�82�0i��m�D�B�L�~�f�kr20HҘ���+|��>� =?aAŔ�mf2w잿U?R7�J���7T_� �3�D׌x����e�%9���ճ���`yJ'u񰼓�"D<vv��OZ�Df���}�B����LZ�Y���P�#!��q5���6뱽Ʋ��mq//���#R��y0Di������$Du�!��|N0?�oF�.k`~AG;�
2�X�*�[Y�j��Y��\�>�X�n��L��9`����'�3׋@�R�>df��40+�^��|ڎ�҄������b�UQ_�<�w:w(��Y
5l5L���k��h�3��W�9s�&�PYH;�LfsAd �	�[�W�l��*0e����H:�gB^�oFa,q����5��b-����\3�߉�ϓ���o��� ó
��������Dz�Ȉ�mk�n���"��o ��\�~�@�M�?'��uު��.+Ku���#�/h"�x�[�'!����U)u��i{-��]9�<JG'b��_�`C��y�l���_�X�ON�CVǨ�=iy��r�s�̈́{��(:���ὴ=��$�@�0*�81q�>����(x㴴�#YhKY{�L���N�P���%�V@h~���ka�d�Й���!�
�
;��-��wn[48�qq��eaWhNBxH���*B�M�4��ҾU�+��^!�����U�(p`�O���@�Γ�5VW=��x�ұ��F�]�:wL� *4�Gɚ���]}`Q�W���,�����v ��`��a�͛
��h�bO]vi�<��rv�u'JȀ[E�Nnlmc�Bk��a�3MtC�?�
�{�K��2X�����PSʗ*�� IM7P\��ɦ�{$��i����}�μ�:?��b���E�Ηx������B��3�`���'.�E ��l����Įb��S��a�NVrTI�;b(Rۚ�3w� O�Cou���sS<�J�Vլ]N1	�����&�-x*!eN��pϪ,?�w�՞�U�t�cѬ˥�JM͑�	CoW|�/o䄀3Q�y��Vsϔ+�H:���c<�؁˰���]^��CJR��‱�]<)�i�*Q8rI]���23�Ċ��L)�{�4U��u�S᱖Fzx�&�**���Cc"�۹��a'9е#X�ࢺ�iA]9��<XZnV�(��'V�v@����i8~X�����y�
��}Ύj��<�M�8-\�|�A֐K�ݑ��B|* ��0I�G*^����J�A�(`��+M��ӎ�.����=X�?b���Q]�;,})�h_��/�o���w�c�i�ɐ����Ԃ�ڨ
�Dg�A���Z�/+���{U�Geo��z��)�H�����3�v{�pG�t�_pna_�����v�D�!x��^9����	��z��[m���b�2�۬7�� %ބ.@&�>��;��3�R�~ʿ`K�xhȦuyke��tPp�e1�`�E{�4~wv8&H^��ˑ�j�R*n<���Sş��hm��8e6�<�Ë�vf>M�f�{��j�E^"	�.�X�$٩Y�c�7���{��n �L%��I���G��S�e�Xi�M4��U�|�L��n8Kņ-�,a�tN�c rg�ytF9\�[] S�$��I$��O)��Q3PWc���	���!qA �� DyTV��*@�o�3v�޽]���{�S��q������L�5��/)�A>$Ӈzv��}Uc�lw��B���k��ܽc�����J�Ź���![n4�g�����qʵ2[A������Y�Xċ�B'�����1�Q�$(�VN �}��ڀm�ÉD�f�[�<.c�'6�����k�=��Y������,ӝ�����`��;4'��8,+�|�b���B��G�8R�V��d��N3؞��	���'�����k8��3D��0˱�N%���[�+���N��Yn��HgLύ9���X�Js����6mnj���n�����J���o��E[R�1����(櫟R(��ɳ�z�v��G7���
�	��E����2m6 ��;4��qć�x�,b�\ڔ�Χ��p��?���v~��[żE��e����H�.
�T�5��O�
?�o�А"��#�nX�@Ҙ�n�~��u���	l��F6ގ����{�0����5#���|�v��E:�&�;�b�C�ܕ�Wi��W�Q7�i�"�D�%�.fJ6:��G�0��-<���~8 �Y
��$�b"FwI����@����vnG)0m�傶��	v"c�-\���i��`�a0�����5f����_r׿�ִ�8�����������`������g�F���߮7c��or��D�>?�%lѴJ�n��K�w���!G�4��ձby��ͼ�G���NnE5 ��6*���g��h��Pb�S����f+�f2j�*t��9�M��M��=���2������I�H��/�Go�NxIc9mۥ^��~>�Ѐ�9�SF�Џ�	�ӥ���@�k�������l�4��R� ���E��X���ԥ���#�c;�����%zQk%_(d�����4�E)��θ�����}\Q�����Ĥȁ@����P�(?BE�N�%e����V��t��i/X�������v�ף'Gt릪/?�B��j��|��=�	k�f�X.LC�T�ؘd�C�.<HY�j�" Z��A�����Zgp�n��Cy�2I��=;��1��x��x\�I� `d�|E8�;C'z�<�O�+;8k~����	#'Pgr$�����SCA��w��ƾɭWb.�R�j��^/XӺ��s�y�DrzL?�1�E���8�,N�[c'L����t�
� i��ݾ�����>Cd �o;��.��7��r���͐3q�Lc�C�����V�1�V��O��<Z`��qϻkI�7����J����8˹��̡<��M��උ<Q�Y�g�K�:4
�Ι�4C�X�M:�X�>EpK�Tk���/�Fh����\I��β���qy�B�����+�2��,$4���W���.�F�+�X��حl�������H:���� �����«�@��X`�y��I�o�o�9詟u)���^rObA���T1f�RK%��=�$��h_�1����h���Q$�V � 4�+rH��ŧ��%�{G���}���r����Թ* Ю���E�ᕼ]4�ś$�`7��"X{W|��D���BSlπ]y�u������o�?��3S��S1\�yʰ��r�[�KN�9��W�r@��8oz*�oH�N1�c���C�2]	nY�+�-��0T_Ș:t݂7IU[:(�#N�tj$�;Ö����B�7xK�#��B�Y�����F����@��d��Q�O��,Ռ���d��K�m��������֣�P�����/��:�(Ws��<\��)`y�|Ź��� �Gf.;�	�r�[���୼�*	 AI�q���-�� ������m��`d�+h��F��X��3ɱ�G�'�Z�4e��CK�1\PE�ȓ�]�$r����%��Ź`�x&2n��	u�5$�$���:�m%a���ge�Ԫ˥"�6�I�o�</���`�!�t�T�^k��|�"a����K{�)?������4��G8V�?�Q�E��IOx���>G��HU�~�x?����1��&�S����e����S��%���C��?ן�Q6S��MhB����L�^d�3 ,�R�Q�%;K�f�q>#�Ȗ�=�� \&��)��|[%����1ϹX����	��;�����O���`U>$�[DIΏ�V{���Xo:t�{�ZԬ�x���0�
�G��O�`R4dݤ�]������k{�dl�hߑ��_Gս���t��-�%��/�j:�b�
����*�A���s�w�?��u�09��k�G�1,��u2���T�m���W�~����!GM�'�^��I�� å���.(��$��Y�N���'C०)$I1���2��p�����luto�!?=΅���িQ/t�U��s)�x�X����>a&&�?����X�`��6��.�[���VM���<�Ѵ�f�To���c�X*��������W�L� �	^��?�Ѭc����	M�Q ��[�����\�?������Z������`�VcN8����C�r{na��En�ʎK�+��Xl�����F�uҊ�[��_\R�eBV���w-��0���j�>f��<��ߡݎ�O�=֩d`g�L�Ih'ល��d�RoD�m�=��? 3�;��@��5��q@����$C\Y؛��l����R"�	���� l�⥑B!?9�f��Y����}���,. ����y|�`	�	%����5�|�rk��L�CZ��0�#v�mpح�-A�6?a"�R��D�U'aK.���)C�gGz���~�/��ʅ֧���9�!���~�N���ȆP��Z�W�1J���U�X��7<����������2͞�'g�?
7{,�?���u���1�Ȅ~�r��� ��������ue�R[�F�ScJ�]}+�Ȓl��oV�I�/|4o"G ����.4H�hM��R/��t�n\3M���ȑ�t'�T�X�X꺗Ģ�xǣ����@�秞��ap}���T>	 h��}��d�`{K���m���_ǰb����d�9]w?<ֻ&y��HH��LS7������uA|�q��!w�!U{t�.���F�}H�6�����_ sϝR6�3[��ԛ�qlT9_+�#>�Bt܈�%ℛ���ɀ���-�Fy�MO?1Z��E�s�Kw�����TZ��wD[�/B	(e�6D��p�	���7&� �����$��E�&�<{pr���\߬v#4[]���	�w����x1�a�0[��Dֲ`8����-�݆E�,x�T�v������ϙ����]	�J����l�;�h�٢[O���\=��@Z}8&O$� �Y͖ꑐ'5F��.�19 �pg��*a0{�;�rh��B`1X3��AFߒ����_�Thez�E~�Rʊh]�u�ġ='��KD�����IUJ�ށ����M�޻�ON�Hꞃ���lU[7#�ϓ��-`.���f=K��Hq>~o�o���ګ������s�)s�m�>%��'=���w)���1�Z��n&���p�h�wC,DP�g\�ؑ�۵1�f��!�<�������	oxI|��e8"|�ٟp�YxzϺ_ZdfK
0�.�<�6B�A�,Ԇ�G�U�����it%��C���#y��,�+�X���� �f *m}��=y��jZ)�9�ml�>B\"�����X�X+�H��M��ّ��:�܅=����E&�N�l짣ߴ��mf~v��M7T2�^A�P\�"�{j��Ŝ9��1f�9	H��ڳ�T���m�[6��:.̇�be�R����~��/�:&��=Hv_̎ڷ]Y�����5���� z%C/����'^c���3;l$�,@�SHD�8��:����y�l��[��F�v!<��<e�0$�3���FgJD�8�9���aP&�P�S��*�,�B�D�$�c�� E�j�� �g`���)z�J���e�<C?#����ohJ�_��E7�;S�u��n�"ҭ�9���F�0�p�Y����7���y���N�'��^���]�������DT �(ҥ���+���qT���y`mg˯�Yj���"2��$��>C��)�Lz�As�� }\F�=F�U��<�T�C�s���o���0_+ݶ,k�?�3���(�FuN��/Ţ�J�%+[�LN�^���_O r	�ʳ��#��C�TXB+I���`�Lii<[���ɑ\���"{v�>A6흇�dpp�j�E�������ˉ�gS�hZ����Ķ?1��,��(�u7�'ep�P�w���/��6y����/�b&^����J�>� �U��x�������R#IFCd��n�)O�T����E�/�Q��7NN�$�uZV�1�uʿ=S]bU�B�CБ�V^��_v�<��T���hk,�>4R��j�L����f-Չ�q��E}�p�56$��^Uz�[�H����æ:ٮ��ˣF�u�V��_�:�?���k�d=w�*M�����Ny�y��L�����>�n�6J���Gp��HG�m3M����\&���,��9� [&��g\d��� X��>� �����ȫ_�����XA�r�L�܆� $ڬ�K5��ᄏ>�u�kJ����iO��&v��#�6�ԌTRڕ$�@�[N�װ�8��*�q�^��y���X�:�@2G&�����C0 ��!��a *�`�\	yl�����^�_��o;7l�fla�2�},����.�T��F�eh�ƮO�D��Ek��+\IVd�%ԋ��!j�]R���&9����$
�#���N�+�G����FT��C���4���A/�z�
66�t�k�i����!� ��ޞ3@p��y6rk?�2	�y�,�²�o����W� �J�1�:^#N�k|���R:��e� d��;��/���(lϳ���ʐ� [#�qR#,��ij�2x$��i��j�a�ȫV�w��Gؐ�%��@V���q��u�b��r�O����nA�C��������,:�|<0C�vɫ�KY+�y���;��+��hI�إc����˃�zB�=��.Ȝ��#|��̜��]��H�ĩ�<��@E��$����s��пf�zc��2=\�_�D��o�s�g���|�� ;���aۢ��d=��
��x�G*���ݷ�
E���[��T0)�8��Fܧ����I��jD��o�)`�]T�݊�R0)�v�"
�a&@h�h��}l=�[��Ӡ1˓���cٙ�&0NGY�\��w��,�kZjZ-��/#a=<�j�p�>���q�h���3��@�&wz@U�r�?�UᖊäW�������:�}t2xT����28��.�[+�Q�S_���#2�����6a��Av^țigyщi܌b�!'P�JzhS�Ϳ�"�B���d~t�c�M���4@��?}��BVh�_h���QPV:ANflvy]��"#5�a�IM��Z��M4�"
�rJ��Vس���/��$�:���u�ZD�C��4����������� �\�}������&�vn��#m�}At��|�(ݵ\�rIaɂdqJ&��b+{��A��%���K���Y%)���b���9�4N�F���yڄ�$�_~L5���{0���^�u�ʹ��?�-�)sm����P�"Buvlp��Ϝ�*�S�P�4r3c��l�S������2�o�5̫�Y��V��c�Ǟ���X�P����h�tw�ΰG�������*�@��q���]k�qo��"TM-�9����s�|WK	��Uc���0�_4��7Ci��5�]9s�8����%4�0&:B����D�(�kd�P|��2 ��$-hl��{c0U5;vA��=r��'�=ߕ���_ː�!��떜O��W	�B<���8��(�׭zd�'e©���i��p�!��7[�������^z��x��D�rVg���hkQ�J�8X*٬�����-����Yc�Q�@�Y�����>�+�"��䨹mvTÏ~�,\��?ݤ�O�AC�`8:�;�ӣc�5%
�;5�i��&<�Q����6u��K%v�Ģw�����}fq�k� �$���;��"�GR+�~<{_e.y���m���yzu����r���+���Iz�����tr̓^�j������S����)� +a��+j��E�:�8/\#���Q���!�έmc� @h���;)ى���zDTĞ���}Ȅ�/�83c~�(�ׂ%g3_�qN"�ե�MH�)��y#��L%�n�A5�aK�J��t'�䬮4���N�+�X��w�wҞ��n�d��&̓rMu}0�"�M
�O�q������r򝾅�������[1C*�>�Q�!� a����j k�QR��0$ݔ���-aK~�HiV�-�%B�B�Ƚ�Ĥ��c�>@�r�ϙ��f@�b�ܤ�ā���E����@�#���'x͘��G�F�p�*��/P�*�}+u�y��!)����	'�����F�1Z��?|��
�VbH�L�M��6��(�@�l�i�
�����hR9�§wf��=��N�<F������w�=�@�0�ʼ��O��^����\J~�('1��	A����I���I0�����NpQ%<g,��:�q��|ob˥w��/�L󚈉��skMI�/���/k+R�&fl�=A**��ܡ�M�g����W4��_���C�в�C������+���<j+[l{��2p���a���:���?��yM2��}��t�������4��O�s���i���=2��Q�n����z�Em��E��G��E��]x1(�_D����]�5ө}m*�~k����5Q½UF��y���ۥ����mT߇yj\�#�5� �����/��Z�!O���>53D�|��2;���m��)Ȝ���u����׆ğ��h����\�Kz��	�j6@�#��R�U j ��ې{Cj���#�{_]n��o ���Ά�\�ڸ���##�Aԏ��4Օ���k�5&�K�5766����	J;P��!���%�TOC�I��{�?Ƕ��g�2{n���Z��&JhJ���s�8��q����9K��p;�pV����/�'Nb\ƹ�Jp7�Ư�fEl/�2�P����b�0Y�O̳`j7�orO�}��R��n?h�Fp�"f��hɻ���a,�����F��Qq�k*��S��~L˾���B�%�n���_�6�d��I�����B2��k6Y~`�`��׵(�D�Á~iX~0� �_La��|E�L���&{�M���	,����%�E��b������!���G5n�Cn�`�TD*�/f�M��W���\ Ц}�9��4hD�Cl�m?�4x�����: �TF��*�A+�2��HN_λ�WtFȝ&����H8�K'���zb�z�xD��~��߭�PL#Bԣ��2Fߢ�����a��"�U�ۨc3e��\"Mށҏ�sG��!B�ˮp������s�a�#�u�G}�x�����_��W�Dj�nh~��b�zv�tX�o`d�%;p�:?7��
��Ѧ/V���|L�Xz�9,�s�@����l����L�E{�*/�X����W�19C[��"�>0�yt:�З�񑤻yld����r"W������J5P�C�7eb[�/Ά�߫(T�'⨁7�I������{�D)�s����FD�N&�ΛbuB,��uW�� �hB{���O8x �����L���Yx�*x�N���C�U����
䏔�yd�lGR�@8�\�e�-w�d@K����K;��DE��`Ī��k������0���>y

�o��Βd'g+M��m�����O��@^ł9b��P�>&a?� ��<�teNU�޶��N͖�թ�r��u�rx#xy���m��D�`�Q�#)n�s�i�+Bb��Z��Iqb���l��<?��5��ɒ�W��.�3����~d�+��ێk��A�͇�d����X,��W��ݽ�=��N�a`7���㽨��#
�%�%,,���`�e^�
��L֞&Ζ�>�J�K�  ���
8�(`}}M��=WVDL���JL3%5���G�����������1�.���ץ�0|��
t�O�����ϛ���-uR�i���HfIqT�(��_X�Y�\����B�1�뉳���J�"�8�\���*��N�8����k�D�2��1�^G�%��^�'2���v9���|�[T��P[��� h�!�*�sZ�
�LN�J���ز�)W�>����͔ɩ%,�Y��}+�J1'6l��4v�ɠ�v��us�sdt�p�9tu��l�X$Va�R���3ګ�"�0�i���a5��`��|ݨ���#Pk�e��[�'>p�
���Y|��gQx�-F�GAǃ}nPN�0�B�Ђ䧩U�PVX��h�Υ�Ռ��%�Ɠ�P�qT�f0F�`(��ye�"���e,œs&�x�����?l��k�㛾2���kj�w���6���Vv��d+� ��_jښ�5Ԓ�2�MO4i�����ڏ��ݷ����ċNb	�M[a�Ft��yo� h�M�ꡆ��(�^���[�]^t�]':-x�_]�[â�[q�ɽ��.�c9��슌�Ǹ��� �p	���28�SG���MLn�Ƣ�Zܐ�����Vg��\�c�v} ��(�^^U��^����!�������K�1�_�0����[,��B�?�-[��h8<�n�|�f�cB�)Y�7'�B)�'���%zY��\�g}x-�u�N�&�R�s�:7
�I.��� tS�N���<5�bl�9T@����x6��t%�b�*o����P!�.I};�������;�62!#Q���y���x����������JH����M�{ٓ�?y?��ȭ��Ə���2c���")�����q��=����Af�}�kY��w��W͏j��3cZ�aWRҺ�7��=�`JSE>`�������4|U&��c��G����ZC�4�`j�5/��g��X�\o�?vw6b�\	'0���}���L��]�
�k����MZ�]�eoF��V�9�I���U"ʋ�cۡ��=�
�x�ɝ]��o	�Ő���h���Y����w��7{��_2������F�v��1��-���݈Q{����3���c!�^�:�r�h�X}�������z�[�^ح|�w����u�	B���X+�[����]a������@R�h.����li�rͫ��r�&�)fW�Q�Q�(�.W�� �CҊ(��i�.���Nď��d�m�<��S:��'�b��Fں(�
���ꢻ�l���ò� ����NO�6EqI_Wl��`���G��!Ǉ�1��C�ֈ��f�|��k��v�gu����5=����z�䥜&����+ʙ��	n
��j���"-n��W�?]��'E"��s�@�] `��~�o^�̗s�;��>��c�2H�jRB�`!:-=.I��xZ��(��0�߿��;�XOb��Ń#�"�5���
�νc�h�+�� P�<�b�9c��ծ*��Sݠ��E���[5i��1`�v�|�м��fr��R�hѺm[{/-�����r��iT�>V�:`&�p�"�G���O�98�U�ח{p�FC.{m���g\�l,=��`2��Qa�U�a:�����*�����di�6jK���&G`ѣT4c��J���GB������s��E��%�����}/��Mv��R�b���+Bٕ��O-T���N�Z??��t{�m�9h��W�u[��T�	���w��9��o�f���aK;G��#�?�bUE�Ԇ��!�}*6D���sl�#��p}.{�&u��ȷ�JD8���� @�1��c������ļx`a��%��ຆl��/g@n>�)�~:���uf=:��Zu5��h�XeY+�}$�9k�F�����C^�o8��-�6��ړ�¨y�yy�?����)&��T-��pp��O��̈I�O���5&�!�E,�cK5�#w��J|9����qd�C�#��Ɗr�h{����B���[�o/d]�<�+IU�=9y���Ζ��r9�h�cM�C��"7^�j��6F�"{��5L��`v�1wS�UL���uM�ñyw� }��B~N�v�mW "QL�H���#+�ĩB»���7�q,���~����W?*��Z�7l��:ƯYLO�%�ǹ����
î����q�ԝ.��q�`�B�)��HY�<�?�N'��z�6�i�1i��U۬56�0L,�{N�Uˏv���:1�F�������� -�M����]���od ��/�I�z�Hp����l��J��j�h1�ރ[# ~�{�J�n���-������TEx�f6�-�\i�dR+V��ׂ�Qʅ��5 ��9F��b�#6HJ�~�[�9x�kȪ�UD�S�m"��O�Gͳ���(7�F6<��c�0	fi�ev�Y�m���f�m������jN�b�n�a9��K6��]�����5�D��pE�L	਺��-j�$m��{�ôܘO�'#7�6v'6��b��ѳH��������"Z�t"�}G��u�C�joiˉ�E(<;�#�/0��ܫ1g���gi,��u��	�n!��Qݺ�E^<P�r]���ۭ/�}\o�U[.i	o4���Ԙ��/X�+�ڳ(�:��SO�7jhu��}��!�![��L�t!�#��؃��l["�q��}P�]�wG��Z4��=X_��x��7V�9�c)����[7������*��dp�<kF��KY��n_5�]<��Á����~�� _�	��R1�rS��%2|B�H'>��4�L��<dd,1���W��)���Ӈ�v-�j$����1�!-�x������t��t���w�(M�	��4D��H�7t*�/�R�:6�u�����&�?���%OF��4������\~Q6mf�tCa9*��]h�����=��_b>�u#2�z��P�������/N�Q�C�]�C�4��_�iZ,��tB��+��bw�V}��Gi�@�Y��'T����/"7݋v�Vm����W?�D1� �$���Z�֋k&��wb�!����A�k�NtSr �75ՠP�M��>�b�|�r ��A	_�r�����U�w�`�@y�z�`Plà �$x��(:J���� ���!���0H�*�3�(�pZ?��j�iG,��Ȣ������q��v�EA�q����D�~�QLq�7_�Kh@�*�H͒�����k�$	�ө� x��N���9��c4:�N�zt;�y�A��0�셪G��O"�۷�-�☑⊯ ��S^4�%�7�����V�],�v��+΃����N0Qp�&�ɍ�|f�P�eLm.�a�a }�,w2�?�%.�@j��[6`{�	E$� �����?��$*tM���Sej��.J��N���������r�ָ�V�q�ą`��k��G����Vx���nj�e�s�۔fBW�@��?>�k0�͡V��1єxGJi�����M����Y��K2��ݾ���>�bR̝]��͛.�J�(�xny�l��Yp�rzۀ26t�CMy�D`�A�����ȁ>Gg©#��E�YX��B�Ome��	�>���s����ߛI�MF�6;0n��o���`��7�H�/i��`�t[fJ��%x�,�K�0��Fn�'��E�L/�5�S��ݕ�C�n�{s`���Ӊ��N��u�!�K�2[�"�lא	��՗��A���6� ��u����m�F�����!��|��צ��To�B=;�
hj7���	G�����/>��	�:��ځq��?4a��o�W9NV٦R`�W�WC7f�x���jo:����� f`�a�u�n�5��L����y>�1�vC��Y���d�������	�k�oE�����X���%�� vJ/ab=5��;����i.Ӕx�0�O<���^&8��	Y�-��$gKA��	�B�%U}v�$�Z��g�1@�y�՚�9�9&�&�RE"]��֤��3����q!>���z���������1��)�=n�V���$:ݻ��'�)��z;�wѨ����<dө�O�,���l����%ɹo7$�ۋM�	�i�N�f��is+��,%�p=x[ ���p���;	>��BW-�=A��j���%���NTA|i�(�B��A�����Ň'���޸��Y��0ٳ�wEmd\�O�<#.��@dۂ+��T���D}o�6�ӄ�ѷ_�~��b��1���4G݋ӌ������[T���C��ܦ��xl�S�Xٍ�y���sYl��d�G � ��C���2u�O%ad��ZV��4"����ԕ�r:4!To�B)}H�3�Q6�'�3�H������f�Jc(�'Jnܛ'��ǆ�i�Y�.��b�%K=ٻTf�q�oʸ��X���sy�/r'�-u�i͗����)���z��֬m�k)&�o)��x؎���g m�+��9���M�W�_CU@���hc )�3���г�k�;��b�.V3Re�\~������̾�nE��}!XjQ�NY�%m0 �Q�i8��!�0�D�co��皵�J�\��׹��*.ЫC��Po8���}���D�lԭq˃z5Io�����K <�C(�����>��̞(ȅ��W-�����������Ax���U�[~�Wj8�ôc'�0��Ƿ97A*��h+�&��jX*��|?8|������nn���%)&l!����7n\������$�(��.E~J�B���dӬ?I�"U��L�˶Qm���z�ksQ���6�b4�셁���9%~�������'������&�HZX�@@�4~�z�T"�|�W%ك�gwT�`���퉷0�h�񢻔Y����{Q�М�bu�W��L��3I�34O�X����܂!���'�t�i�Q�I��������bӢ��E��u�J^���W��E(ӛ(]�J��	���c��-���}�@Q�L��b�����{���b[�*����mλmC��Z"��6�4�Ve��;f�'�|h���ג[/ͤ ht�o�/%)�]��v S�߲������'tԍjܼ���&&�����ۿ���Q$TF���!N���m���b�@c� 2��h+����XJ���9��j-@���	2t�G��^�:���?��2��،����"�h��p������C��g�n����(>*��#d�]�v�>)����\D�͈��Ir�-sξ�y���$EL�������h�������o����sd���+%d[q��n5�\�<˂{�J֊2@��)[�Wp�tT��=ʮ��D/3��'%��-l�}��Q����č�'-GU�Wk�Z��|�|N c�X��k�|S��)T�Iz�D��E�I������Z|rl#¥��ݢK��M�>��I�CmF�#i�.0Q�2O���y������hp.��tZ�t&���*����MY��l���''��:2��{F05�b�~Ŧ��٫�u������y��\��;MI��]�(~r���w���A���Y�"�3�>j��$Hd5.�+�4�ы��3��!<[~�vȳ�R�^P"Y�	%�AQaW�ܸS�}�G��m;�8JQ�@<��Ԑ�0z�Q������ܻx���=��g����P�w�6LX�}k�����K�
��r��l*ꅟ�3(��B�e. ���v$rȸT�	�_�\�'��F�j�ܢL1��y竂�ա�����.f�~�����:6On�p�����br��1��	��(�0�I�`]�`N����9w ́���W��0�,y޽�9�G��qv-s�i�b�1����::�\=�l��t�2oڗ��׊�r���.��ȿ���P����fN2�o:>DrHߕ}� �Vi�y�jQ.���i��Q���õB��T�2��l�1�`���������aSmP�OW@��Mf����r�8O��X�
	���B�U�c�����$Yxc���剔O`����'H."#v�5�g����=F�	��Õ�a��t}i�I!	�kF|�����ǰ�~��N��<����%ہ�(2n�M�v_�<zdn()�۹�~F&�CGL����f:Pxt7<ݣ�����Q/�5�<�ˬYF*��5J��	f��A�V}�..���Vp���y	���с ��U�\.r;dga̺���tQ���C4r*H��}����c�:�׷��!~��e�� �J�Mv #?�����.~�9^,����³c������7V!O�Bn-��0�Z��;d���v�&�hk��N�\���'��N:$��%#:�Ǆ������/u��"x��۾kr5�&3*Vo�������%$a�I�G���SA,��CD&��,�ÕGn)�%R�q�Cf���^Q��z!껶���O����r��*A��k���2O�Lh�l�0�Nt�h�w#W?x��;�(]���A���q�dw)3вh�6�/?��a]G[�V�3u���]��'�?�����hMrF�,}=������y�i:�D���dr�S����Ia�)pHV;�QB'�W]p���P�:��y�7�qEpb6������wxm��͐s�:WJ%�V	�_�Չ�'���l����ޕz�P�B���<�[&ݭ���H��yL�\�
걟��9��Ys�L�n�ƶ�6t�j���L�B���aF��3��=�Fz��
m�7�DA�J��������q�cSkSmA���(��aȮd�(�ք[A������B5kj?*���Ub(���U[�n��G/*9����$O���D���h~�|�+�ȯx�`+l|f����I#�5Do��j/�v��,�	l�YYR}/�>C�kn~|����<��>�	�_��{,W�a�w�U�1�&�k)(��f�I~��d�4�<`oRwm_�����|��v�*��}�j�-�g-(�۠� 	���j-%��WT�o aM<O ��K��ȝ1a��:�����jõ`d���v��!�efwf��αk�	�:��-S;��@�E�KX�qVRt=wz�O��yk�f����<n@<�4�>�S���ެVo\�}d���r5�<�c�����ب�#��!#�$���1H�J�p��hcq��_����C�9���$	ʁ!�R�"�]6���`��UU~ak��Ƌ�e+B�WE­u�Xd�	Y%Uy�,�3>�-&�S���xs��?�i�jR�� �;'�F��ئR.����)�D��ɕ9�}^�C�-�s�j_;#+H�;Ѵ�%z�q����ˊK��B����k�ڟ*Jp
V*V�s�P�w��b�XW�3�Ǝ��H�Ӡ����@�D�ʬh�iQ^0���7����? ->�G>E{v���Zռ�i�&
��p���������������ϰ_^��5�p��m#�E:2u���ਬQX{�K5�#u
��7bWN�A�40ᣓ������LI�猼�n-B���� ���{&�ޮ#P���d{���Hj�*�N6U���H��{�d& yܱT����(���*x� �<M,�;�/��+���g"Xͤ�?�dШ�`�mdgڰ�V.^�u�t1�0�H=0�w4��n������o˰���e� ��K���b���n����7�&G�>ԗ-�;ʰ��E槓�������K��V�f~�0K��;/Xf<� 1�1{�[�;Sg��/;�a�}��nqu�NC,-0�F^	Ӆec���db?�OjVl���m�q)ƣj�Kb��_y�m� �8��c���?��R��t=��7�r-8�O���`��V|��e�+�]��y�5T���dԛ"�o��d6�Ɣ�����AK��S���������$��} 3��C1�HΌ��>&,�`��6V�_�:��f?�;�B!��@.6�cX��]㪴��}%..ir^�\v&�戔��w�V�����;	Ws�P[i�����O>ַ\�?�.F�Rck���������ȑ-4,�P�Y>=w�e�i����$��I:ZSy��ZR)m^Bo�|��-�S��,?��G2U;�o��h�愛�#b��h.,�aq��W7Fj0�q�CA�C���A��(��d��_�a���.g����w�P��u��YU9��\ޡP�,L�����OÜ��!H����"̴@Ȥ<�hKJ�R����o��O�[Wi��o#�fu���#��9ge?M��׋���h���o�4s���=`il��Z�
���>������f\��g����Ͳ�G��F������o�U�7	�����l_���ɸ`����@V
����LyQ6�����d��V�|����h�f�8�v2��+3fv�VL� ��mY\=�k�vj<J��xg��(�I��lpNVU�ę���������̎�PM1+�4	[�����}�{��!��Q+���v��|?Gp�ކ����b.4;`;�o�g)g�4�(GX�Z!w��P=����'Yn�m_����>�nW�* W�wV��t@���ZD�G�&
��Ճ��R�<��03� ZOI�Ppk��y���`-����g�]����:E`��5�}����\�����L�C�#��YdaY|�&T.#��8��p�����*X�Qs߽��K}3b5���GF�P2�ѿR�F�*	\=����'��ȝ��"����S��\x|������IN��
8�.�|�o���/W���F�\���?g��ric���1\�~�I�Z�Y��~�w�|t(�9�$�к�H�hp�(J��k	�I���?�lLX�O��\Y����=�d�;�oŸd^�]�~4�&p�V����`���wu�%���|� �Xf%�x��I�K�����z���x��.,!����-W^'~�ۑ���>�=<=�As��:�V����~�ƿVJ�n�C���L����>ב�)]aH�I(�*S[B�5�2����ޙ1h�m<\�:f�[�3;= ���.;ɯ��~-FAN�P�U��v��h��/ϰl�1�US!�gy�s�5:�����8�W/q����4�ę�bƠ�hU�|�=��+���s؅ �TD�_FU��%H�f2>�;F'1��C3n:�a�Row��$vI����������%L��eY���B�.�/a���v����<א}�~�˨���?��:Qt
7H��Q3���
�/-��Ý�V�u؆۟M3M��f`��)=�&X����*�	g�Py��yN�q	�4�blҁ�ˎ�WR5�u,���ً1�}r�F:'�C3�#�f�p7c�Kժs:��O���T�k��d��k�#T�|Dl|��GDj7X�KU�;�'6 +���=��n[ w��a���b��O��U��=©.,YH ���.X��s�z'I��3���4Ib�鯨�lA�;1�1�f���%Ux�>v�⻙#|$(����Ј�	b�wd4�D�����]����gU+��+���x�ŪK+�/��7hu���&+��^@bU�R.@��s��9;�T4�kQ�U밆k�a�B�z���J߄`�U�0��.y}��>s6����_��Yq�b��6Zr�9�������}�j�sVwb^
���on���a���9�KY�q�A���z7�h	�]b�.�~�]C�9\�����ыíp>:��r�}}�7x �W���nxY!$�8z��~��鿲Qʈ;3B���3�P�/���g��u��^��&oS$3�ʐ�iT�_����B��
-,�a��w!n������@hT�Ms�z"ޯ_�3�n��=U(���4w;j�fu��X��� �}%�u�*��}7�-�������y���}j���:����$k:τ�σ��ٶp尘Ѕ�
���x��mMH�4Q���ڊ���I��3���T�J�t	� �T�2�׽>�k|�0�Q��h~C�
�����N��� 6#��]�x��JiW^��Q�7S��@0�� T4
G!��|2��M�B�?�Pq:%�O���������z�[1��U6#�2܌�uħ����Z����V�z�s� ������ ���e{�gC�+|�w�$U<�2 �7�������8�t�Ž(N�Cʫ�m1<�e�Te��}5�K
�����@�*��#��t��i��Wu'�[���vi 	`�ڟ�9��]�sȳ��rz�H�3�j�pKǗ��(X3���D'̼g��$a]p�v�ܘ�=�ׅ�]P�H�;b�i'���~؀CY���Q�Zߜ��X�}3��;�%�ة�C I^���o�lB���'ێù�#�����1T���l쑥x[��$��\L2v
�Gh�-x������ �X��@�4)�Z~a�!b�fS��B|y��|����W^�2�V�.u�Ȁ�g�M�J�*�³�~7���[�q��_U�Ց��f53�;fX��l�����o��˩���4ԕr�ϋ�	g(�����nRh>�q1M�ђ��Z�A���G�Y,2���Pl懖S���݇�#�]� `Kn���\�[ jy4�r�����Q�l�@]I;J�h��<Y��������_�_$�)5�8�5�g�Y�,ϼ�JuB���*vװw�����ɡ4z6N$;n��W�(�G�fgG�g���8�{�����)�q8�P���7��9����]����܊D}yo��?x�JX�6���s�&:�'/�tۋ���!F�;���'���`75MQ�A��30\ά'���bPxT�䧦��R6�Y�cPk�;d������W�r�U@���[�!����f�e�s�@V3������n�J{���U��6{v-:~�jR���P�X.X]�]�r���"�)"�F�_�Hy����w?
��k�ǥ�;��e��hH�T��v�ֆ֫�D�$)Яe�8i��y���^���&-?��s�*.)�m>-���0��_����"U9�av�<Tī�nV�o~S��à��Uw$o�a!�!ڗ@���Xm�XX�8B�A��p��dO�H� 8G��K�ב3+e�ĩ����p"���OQ���
�WYaf�ӄ�c!�_$��%fؽ��h������i�������0�(�I6'�&Y�w<�����J)�U�e���
��/	F��?�Z���J	��W�tG����ŧ���"�9 ��?�G@$ht6��Ϟģ�c�}_	���'f��	c��.6���׿+�(YJ����"�	�E}?��� G�u[υP��f�F��v3G��ׇ�w��+�. L1 W��L��-�t�i!�b5�lɣ�q �El	8�}BD�h��,A��A��J��O������9��T��w\8�g�{��naI�F��/�������䶁�l��PI�����������Ζ�7C�'X�7N7B��{�.>]�n��$k;�wfz�đ}(����J�(�j5�a#�|q�Ж�c8]Nk�}�I�e� p۵�O9 ?v)b[t���b��J�e�C��2�i���?<�+���������p .��TVZ��n	���=�O�Q���߸���G �@���#��2�dt"����>��ϛ%$��\��4x��}eH�8�L��q��A��7|ޠ�L"��^vsz ���i��Q�OKz;\�Q��ޤ��
����9ZqR�/��"p@w�'��PuǏv�6�b,�T��G�'jJ��Ƈ��<x��,�k)z��S��b�p1��d��(׸����r��IXտ�L}`�]�,~��� �}G���N�vz]���v�mb44��c�{�y�ஈ>�I��J��ݯH���m�[b���2��C��5����Z��h��y,p\�Vu#f�(;猹�X��y\J~��*��*b�|�?^��U{g��ZqV-Y; ��M�����)V�Ҟ�-V�IRh[�y�sM���1s~VDvѲm�#���^��C�����q5E����٤#��z��i E'ͪ�
�z��gjO�dW�����3=7�x6Z�m�N���r�J�B��S�4{�	�,�%�F+G�еy�/�ǢF��ߺ�U�U�=��d����JC�S��N�ϐ��I�6S?*2۷�ޮ��"�9v^�=>�~"e9],2N`ȁv�[c�) XF��"YM�f(�a���$�?��R�(���i������i�kb���l��T�}D:�Q���7�M3$v��$��}uvY��Qqmo#S7}dJʳ�U�E�M�bw<Rbx��˕��p���:L�6�����')�S�����]_�}�ݽ\\�܌��_\��]�o8B�dU�����H�S)�=�]���g����Wܽ8��a\�w����5�tw�Ev.���1B�7���H�_����Ud��$*X3��c��������tډ���D=�1�Qnx�rs�s���q�-����Z�ϗm�zz��l`�J�.*�6���,�t$�J���H�w�.j+�y�Լ�]DO���
�f����2 >��7���(^�3M�*,#?��"��Xv>/˴���<�-=Ol�y�^~o��F��4�*7�)�E���T%և���h�=]���r�9��.U��w5�Ú8�Nh��3Pf�N�_ +�A��,~�@�1ng�ǰLn0I�*7b!��ѥ�ߵ��z<W�;�_��'��4Z�T�mZ��a�O�tӭ!���c0"�]o1��d=��**���4��_��[��"~���F��{;�2���3"
$������P�w�$;"y�~4 ��%�EG<���RV��q݀�8cx@VA��+Y��+i*D�^8�X#ی=O�da��|�����?���-#�|���|w���^H�ް�׍\�UA�Sݟ��!�B�Dy��v�
� ߆/[��1r�֟N�w�� W�Y�`St�V�4~~!%� R]ɛ�_��e��n#Ϋ�%ݖ9�-Y���0�����E)k������H�e�,A��ǅ�}�~#�zKr�����F�x��'�E�-%����`圹J�Y���M��ؿ�g5հ�)'�]����?�v�_p��R4g �-Ӂi�%E좫TSe͒�š�� ���Si��Kw����{��M=��8Gt�$K�=�?@��0L�a����{p~>;���tǥ��b�
�Ϝ�݅�j�R�E�e�_ҬB��h�,�<7@�b��\Q�S��X���9V��˒dSu��fP��"Na�����H'&�V�L�ܟ����p��b��ܔ�fBd�rB�8w�����M�,N�?Z:���UI	���R!�l�7)]�/cw���)݅��R%ų�k;]�,�3�͟[��yAK��i����M�$s��~�җ��D��T3/��`X"Dy2=���QC!6��%����٭�v�1���bV�˟��w�$�氤#����c�:��>�!"���f�d9է�F0��P,��Ra���+�Y+zI�B|�>����+ 3�pfNfU�n�,��� ���7���>�6��S8'H`|�ެv�M����jF� ��@���Ã��Sm�aj�����(���?���Z�v�#zZ�`������|�����L�3[��7��X�l���|�a��a$N�Q���,�e��=:3"���n����R��.��LF�Ay���D�&�s�Ǭ`wS� ��:*�*Fi� e��
�\,U3^��VO.%!J��p[���̏�\b�X�����>�����,�R�L2�����i6�4�M�˻j��	��!-�B�k猷�o߹�P�TU�2o��Z�g +��@ �R�ʹa��W���:؃߽�g�pmS�@
��]d{��'���.�LG����"���X��\��	x�L��.��J�1\]h�#3�V�6y��J8w��dJ�i=K
`AΓ��G��G$����bX.׋<1���~i� �&�<��xβK�&,mU;���o�2*�n��qa��EF��5�L~o�R�^g�H�@�/Q#�ɸ!}���cwY��>d�}蕮�$U�N�q>F�V���1\	x�@z �7�]g�l?�ͭ2k/�����F�i��(͜tP~l�S7_c)@C�^����:��YvA/1���G�*r=�Ii2�Z3,T�=��͐��g��~�at���Z�����4tTb��qm��B�$/ԏ�*P�� ��KuC2-����O!�U2��@oz��*������!B���%0�5��~��w�,�.�4k�0�@�ۼ�Ga X�a�*P���������t���� �������s|�q��C$9(j��j�%�b���5�ѳ��dZ���ܪW9�[:V&*��	eh�PhX��;x`��o~��i���&�%͌>� J���h���QDR���O�R��,/S4�d3��/����v���İ�7��d�R� T%O�d���*��gW�X�{h��=z��X�7��%����WWZ6m:��a��--�{��͒t���'S�J���m���֣!�a]a������qY �0?^j�B���p3g>{|�y.��,_ �u�qʤ��ZzK�A� �~�G�fq�f�j��u�7���b[{�+��g0�~>ܤ���d� s/��
�` ��Y�N��] �fj �,��,�/3P�a���L'Oʇ_]�U�s���ԉ ��lwH��?[��I�e>}C�(7�����P�H�.)_����v� ����-?�"�(4d��L%�,���;}c���}p�m݂�s�
Ct�	��H���<][���m 	��F���(*���Z+� ��X+	;��u��Z!��$o8f�ߓ�S��̸�x	c녻���5	xI��!�৽�~�Q[rx����@m��@�z�n�!%-/�.����<���_�+����P*?�+�  o���K�����x����GN�u����j\���I�&��7��i#�wC�S����Iݨ�Kͪ�f%��|��\夽v��k�
�T���a��Bp6'7!e�/�x784� S� ��Mz��_��䃙�a㙆�s	��Z+����U���lD��PB�Ԇ+3��Z�����[+�Y�E!~��#,����@Z|E��rm��]a=��2>��Q%�(3��>g�hDp��6O ~��ƣ�u �� �|%f	f�9�S�4w��|bo���	D���ۖ�"hqhF]��m��)E`��u&>[Ȇ�qWf���q"м��߂�g�P�����נ�_B��
���lޒ
#�)�cS��\L!��x�r;�������ɣ߂T]�9A�Fϐ�wЦ���+ۂ�Ư��X��/ۄ�T-�e��ܤ�D�9����QX���
��Ļ"�k�k��/�ϖbZ[P^���p��/��QCc5b��|��+J���C؁P�~�K������R"uq����Y�(P�%��&��G�8]	K�W�ҟ}1��-g��r�Pn�'�߿F�����g�Č��ŰÄ�RDrN�6䳙��Zd5��\����e�C�墍��Xr���r#`��Q�������!�߸n��~�b(�]���p�c�w)�ƢX�2.b1��?����#�fŘ�ވ��%�gR'�C?Pv4(��`�)�+���g3�T�n�X�dD��Ny6�G��Z�'�(0({�:\)Y�o<䚝W{�ҁ �^�͝T#��W@�l$���y�_�V=�g�etF�!&�ahY�S �Q��G��7� "�M�lif���H(��!lQ6$VA{3OgV��k1Y��0�0����\1A�|K��#�����4����p�_QЇ.�{Ȝ)��/C{cj�f'�����b�%Kk����k��\~��
��?B8�[��N��$;�_4�+�4:�|����^�uݢ�5.��2�$&��
��� �0�o݋A��ˁ_`�i�����M��cO��1b9�4P��؊�>����n�R+R�L���O`�u�w�]K����g_Wd$ڈ���B?���I�&_�7��r�,X�]�
��B���<3|*/[1��V>Jx0Gf��#�mxKo]ȋ�v��=����AҮ4'�9_SEbm&�^������J�Π����o�,/��im��%�ʖ21�d܏6�D���AV� �{J�6�D��Fhvn��"ޠ�������¿���(h}����G�k�mq��s�Y�x����	@_�`&RR�4����n�y{�k.W7��g����VxV��T�+���je�c,��׍��#Y�r��H��!�-c~�������ߚ�<�\6#�Pw�\����C�arP�%�;���7�@��AM<G^���߅�K�o�hZ�ʥݧ_��W�0n�I�a"~&����%�Z	�8q�A�%J��E�A�3� ��f!̟U�T{�H��L�+�8(ic�"��ܵ��ӱ��|�G:c�-<l!�����0�v�*Pw�Z-մ�۶)2 �0�ń���r
�n(m�]�����4S��N M���fl����r�xf�!Z���`n��l7-:����L�T�bw�^]. �DmwPf�%��.��5��Av�^uh��z���S�r9;��0B�ڮ�3]�����{?�S�*��P���v��]s�����ŭ�А��ڗ����`�;!�ev%��{]���ܡ�3h�y9��	�k�`գ�`��V""��M'�^�Xy�O�I���=����پ����&�Y�z��>f�5k�
�ŷA��{�ę�.m_=���ӗ��٥��~�(��������c�%l@J7���`��!�b>��!r��sXS���&�n�h��\�צ�a�M��1�
�/�tY[�;��r��Tg�ȇV�����FW��+�W�Q�;1��hY|������c���\e�`�4_ČW�Y;M�Z��h��?��B�vB�S�X�A�`�/��HG dۨ��RÚM�`&��J>bPD�8�S6S�C �)�wx�/���no�ʭ�x�.�ɡ��1j�eˀZ�>��Xw*�m�4�>W�%>����䑠r��_����{��D�.\�&���{��u���㽕A{��E���f��%X�%7i�����),t0�:��")��U#%�u��J�cd=��+	�Ǻ���8�@���R���9]R>�A�����~�& ��-PF���c����
�0�e3��h�q� ľ����ʚ�G��@nF��=�Ep���t{dE��_5w��n�<~z��&<��\V0��,m@���	Mh"��8d�/��"��Nl���VrS��I=d_�ˤl�w�q�Aq���B�'�R-Kàp��p��ϡ/�|�����&���_S�u�$�`Nat����R�+�9��d�9<���4.~�ؒ�R(��{k��jl#NF�& ��9b���F���W�s��b�9^��:bɞ_]��D�3Lg�V�)1�'��c���������UJlJD��ƧO�����'��V
��e���kW_}����5ׯu��A|%h��������y`##�q1@�����Ip�Ś/_�*��c��'+����P"���`뽞�Z@�gO;̏�*L��\*��.��m�y�'du���v�܎�ƀk��X���;�/��(���f�f V�1\�P�k9@��`�����_Flnf��E?����v)�'�Q&�UQgR��x{#���.}*+�����㼂�����m�j���;�JS�:XJh� �? /�r/XԵ�ɕ�Q��k4�j�~���3��7�&�bw�S�z<J���29��F?x�}�|^UpD;p�����$�ƹ�a,�ᭁ���㪁��i_I��M��G��R�#��u��g�A�����������kY��S���U��*�J��R!�NO�@h4�ڡ��rZ|.`-�(�Z(�!�,�$t�I%���y���dE��ۓVe��۩�
'VH����f�X�WD�:�[�u��g�Ww��E��� ��؅�jk��~.O��;��̙!�5E��I��+���:�'3�*�U~�m?@f2	4+�m��)���c
�B]�<���=n=�'����
 p�(�6)F����`y���K�N!)��!�'��bm�v+�!��bm��O�4*�%�x�p��W/�>�c���km��\�?��8 ����|6��aV;j*��1��c��|Z��ŧ���z >��7nMG��P�A�:hz��X�H����G荦w#�2���>���,'ؙ!���e:Xg�V)��$v2ÿ�М*ho@J]�Z����\�@�o��f>\��HW�{��"�_�OPKwk�|(�	���|+��_�\�3�N�[�̓�_R_!��C���Z��υ^���,�Y�A
/� j�����zs�֐1Di��T�@4&�g�ZC/]$�:� ���?5J�}ڋZ@-���3ra#Ӳ-���QW����ys�k�mH���vKr+[ܰ�,����ᕢ1�1��?J�+v#�6��'�P�a��Yl��?^.�f.��	H&��P�1:��a���_�_��2�f�	���.��	��"��� �Q9)����Zd�a�0�P4��wC���9����޳Y>+F����Įmd�xS��xey�j-Ǥ�#��<�$�n).TaT �>��S�*���|�w�ZY�M�mK���w!�ܾ"
�y<�������/7V8M2��i�^�ș5Y�G�/�Y�z	�,��U��㯰�\
X� !�gJӽ�*C�*��U��$,��e��_��j�Sxӭ �L`��f�N���(���4kߜ�64�EB>���W�6m�'���.p?���
�z�Oc����o>�P�Y�c{�oթ���һ�E�P b�&�=>����/��-+��JIN�M
B��~_nԔ۷0�n��艅پ��6�/�ڄi(��*���n����Sx^�| 壭�����g���?;�95,O2(u���,�b>��e���V�G�W?r�9��{Ы9�ϋB��u{�1j�Ǩ�G)X���yP(��p�����l`t^�N���{o�S���ƚ��Y�Hڰ�_�V,�[=�u���ki�E>�����0� �q@�)�D�ƥ*��n	��.�A�V>��	��׈@����B�̇��Ƹj�O�I���V=�e|k���=�-�?��O@�"�(i���W�Ve�Xd�$�04G���a"媑�g�z<���Ų��x�Lb����9Tf��`�N����P�ӿvP��u�7) F6��[gx�8M:�H�!��iUhc������N���ɢk�ǡ�u���ǿ?e��+L��9�����-7���<�V�пI4�܈"yD�Y;�n3p�����)A
�+��[������N��u����oV�Q~�v;bZr5�
�׳��A�	i���"�ŎJo�>��z�|h@&�����G'�ˢ�1��6����j0^��Vqq��g�2�$��
�Gsh~���-�_�[!�Ʋ��߹���;����Վ6��m	q7��aY��b��9�X�oY�H�ɚ��SjȪ\����l�p<ژV�c��Q_�uU9��c�֫�i��;��I�Њ��b�[Ix�;���ō(��e�E��µ�a���9���D�Z80$���{Ά��u/�l<��<��лBD/.�T(�M���'��  J'w�䚵��[�/Y�}3i�$�qeC��L�LE%�����b��Q�5���9�[6l�Z6
��n��1�y��l�yr�x�Qh�9�I:c�پ
حE�iF���HLH�_�oX�����[RH�FcP�?l��W?`�8�3�G���mc�3"}<�C���ڡE��6��-������:ff���Gy
I�>����F�F�%�O��XY��ũfPM�Q��bD��{��D쿪�u�4�
H/��G�_�V~����H��m���4�@m�<��h^x+���1-5���i\��~>vM���7��|�6(jZM
�z@�q���@ ����}Dr���l����������X��Ͽ��$�ծ�})RX�v����F��\�����H��T�Qz8��~>ú{J�L�9SpW�u�#�؋�ӌ��������������w|�����6�ǻch��<-jvz@�ʯ���,]I<�Gt%�_��G,����-�/G�cE���,
{G]�%��u'rJ:�Ǌ���R�g��!�7�b5�����V-=3ݍ�w���!yh����<���u�Q�d�52�P޶@�Z��
paOߺq�"Ww�?Gc@]LHY��F�D�c�Z��7:�ڃ�	����C'[0�r�.����>/���(U�T'V�{�f�2����x�^K,�f�]$0����M.u�c���/k��hf��>�8����N	� ����'I��dy�1R&�\��v�R.��U��XC��S�@��HCp��]�(��gK�[LZCD;�r�S��\���h���q׃\+*L ���,�w��5�y�$�ۘ�磔�s��3n-��߄��]d�Y�����Dy�MԖ	�3��49���.�0�`s'����j�Y��b���^��h�v)D�����E~��	K)������������4��;��W��z�e}xr�+�6o��Ɲ��hzX�b�_��D΄�?�yE��������u�a���@@�|�N��M���&".~<�K𱶂�d�>�NT}Τ��+�cp >�ϐ�H
wQ���ir��mk�TN�b�/��k���/�NB�9-2FM3�{IX�/�H����8��u����Y,�Y���c��ɒPJ/�z^��0Ҳ�%K6��K��=��>��c��<x9�܍��(�mR�.JȀs�Ȣ���C�R}	����	lY�z��� ͂X�b�u�IWr�9�n�E�ρY�D\+I�n,T��xw1��EC?��� ��y�3N��)ɒY�Kut�WxO�Q�jKÐ�︷� y�.� .q=�cO\]�Ω�C�4'����+�u�W.^��a���z6�����O�2o������)��
�x�# /#ӏ��\)�����?���^k�L�w�*�Cȉq�q���V�C�;���v�|�o!�����H*�Aύ�0vVi/FH�.��e߷J �O��5�H�1����r������Fn�ù ~�W��-1����.�U�7��	��绷�M�Vi6x��]�:E[?�t8��YR��
��Yn[w��a��a�#�r��r���u�� vWR$�~��������{�����j]X?K����D�$��n�h?���9l�
��󔷯eXC�}g-��u ��̎ZЯoU0�ݯb�H?�&����� #�"W\��p3!%c��r^l~r���3�Xⷑ��:�7�����w��2lM��N���i�UaOr;�An0���s{�
0�!��<e5CZ\z���D�f����vP�01�p~9�T|��k�� [�{���G�Zf���1�z_g�P����R��s�I�`4�27����ʩV�圉>�C��(�|��T�5�lc� C�so�q�uen�g6��6ؑc�/����/�{T����	�@s��)��A ��z�73AHR�$���o~�(~g��B���,��ޜB���8����:��j���b%x���"��Q��w���)n)��U]+Yмe�	/�߅	��x�y(�Mo-M���6�<ެ[|�\���Lt�d�_�>2+L:��B7���q�)�f������+> �@�%ON�g&�q�Io)�X��FUv����2�:F�t%je9��P;{�no�����/��hJ�Wz�7���p�F���唖%���F�����َb/7� pvU
���L�$�0�1W�jd`�8�qP�P��um���fq-�>F�ܽ����"(P{�29q�u�[Iv;Ͽy�Ғ&��f�g�P��/I�!1��x���XL�Ŭ[z��	'��xn��J��[dnq����衣��'�b�~��U��l�{Ć�������r�:�#�,�@+봴������%�,xVj=�����WtE3c�s}-6��u�鰽�hN��q�_�u?�T�E�\D0���kH�fnG
���v4�8�"���U����9����#���wc]q��h��j�7�2qd;%l�jY��l�X>�6t�������0�	�+>�J�����Q�2����Ai���7qT��.���%@$(�zhف��#W�_G��٣[��-�d�sg/@L�!���Q�Ԋ�1xم�o�53KYCr�Fr15T�l!6t��� ¿�i�[��9�w&1_4U�#�����B�q/q��R����톜�3ˆ{\;�kV��vs��.�f��S߫ieGWE��_�S�`�HKeZ�Y�]��K���ccz𽡮88��:3�Y%8���O�-��v�/�0<��%�dF�?���[���FEX��"B�,���"^"��Ɩqh�[�~(���
��T�
����Wf���#=�"�Mh�Lk�$;"&��6$�P��f�MAՎ*�nOlvɠ�+��	<kq�e��c��G&Џw=o�P��,ce�\����g�,y=����ַ��մ��;"Ko���R��糐�x��
{���&�q6L�OP#�hX�R��h������-'�C(^U�@K��?���"=��t��0�b5��(F�et�����
���e�y�!���z23:#�iGn^��^�gC��9�3j�ĵ\ŋ�Ԓx��,��7��1Tok!���d�$���O
�#��$��o%�}� �.��tVy� �!�/"���R�C�ƚ;荫�T��s��j��d�d�Ż��=�s�[�ȸ��4Ȓf��JB���ݥ(����Y�1 �H�zv�v�x��P��?�&��%�@o�-ƨ�	H[&"q{�.�L{���c
S�A���/�`�xA%�&(����4vր:��ev�r�t�D(E�XA���;�I?S,B�0��F�4{1��5��ϲ��r���Anb��H5l8O�� ��YXkTgV�}KiBE�N�2��+�����7T��pj�h���d�k|����js&J��eQ�1f�yϹ
nݡMhg%^�ɠ�u7�;�&��8Z��SC!S��Ȯ|��^��K����ESu����I٩ AβIY*��a3��#"0O�*�G;�����Gن�|O7�����w�H��ďt9x;���T�r;�4��Td������W*U��ߤ��v
5���� k7�PǡԂK�����"��`�;n"����d����U���)R�k�	�5!�,Z��OCZ�FY�j}^�v�΀�n�Y�#ET-������w R�-Y���l0w�T��{Y�����/�=����Y�i*Wf`S(�U�\d����v���g!�$��ߗ��Vב��I.1l�$-m���`QZRg��z�m�pwսYL�1)�h�|����?O�"�U�f��9V��x.m�C �����l��|�<2I����j��JQk�'�� tZ�9�f��ľ������w�	G��qܐ�FH�ڏ���;p�-J#���:{��"-���ӏ�+K�Z�7��5�GӤ��sЂ�����*��]N�u�`P�d'):�U�p�l��mf��jw)&�(إH˃��7ƊR�`Q�x�j5��[G���I=���[�KQ��oJe0Ȅ������IK�l��t�u%���Y��z�����s���p�-�A<Ȏ�I/��x�������.���kA��-c�̪ݡzOH*�qZ��e�kԯ-/��h���C��!T�S��$0�n]���_���1''n�,��y�E@�3{Ӳ�� ]�r�l|�])�=�ޑ���q�x��3��P��`d２2����z�3�}3�U���0X@^���
5Y{�%~��޸�$��[-�p��tܷ��J��i�tlF5J��bjޗ�Ðm��V�Q t����#1'��<���K9U6xqۍ0�|;fei0�s�ē#�����| ]BuۍO_�Zo��=c��^=r��������n�<��ߌ�?�Y����pr:%7jH&�X%�>����q��\�岆�O��Ut*�[�� h�;�.��#H.�ߵ��fڍx�'�묁
O��BU\j�p��ɣ.�Ⱥ��r�4�����fT�,������[�%pC<�K��A�]��I���=:����@��� ����Y��ddU�ߍ�۩&9B����F`o��<^,r��]�ޒy��p3#j��M*jE��_��~����;|��y#�jFb�\��U>����T��[�z+��xz%[��L:���eY�?&���$8,��E�$5M.��aFs�y���i�����P�ȝP&�$*S��;�킛}]w��d]]�A���=�9�k�U���U���8�\>���j����7.7��B,��$X��S��F}�j��tri W�,�b��`9��kD�������^C��q"�M��f�>�yL��J�	 l�\��^��!:�/�_��ӹ���6�����Jm<����1c!,�X��z���/��F��<Ծ>I�*'�!��Ra͛���z ��8F� ��~�D�n�$�ecD�=v��
Ll�U65B�.8g�u��Ǐ��du�|y�<�.�~j���6�,�q<��=�A�QU�g��	���P	��2�����
���3ׁ-ѧ���_��GQ?ѦW뱙��[����2�(��X+�5��V��m�Nw�D�M�kx�0�'/d�C����D�|m��?��hÅ^��-������S��\�m�Q��`;DJ�`���`\1#���,��UC��6,�ʞ"Jw�!���c��]S���Re@��3��7�E����n�\G��)"#Ak6��x��/;��<l9y7P&ly$�;7X7:8��>��|��)
?Q���%�0'�n��.�Qq��\Ȍ����|(�]G�T>�� �R_��Tw�f�T=#���̲Đ�x��ec����G����J$�w�ˀd�y`�S�������:W�&��a�n6x�q�8}�2�l7�/�B>fPYnVx���gDQ&��)�e�0V]�3�ZI��.�Q*�y�jPb;c��<��y���_nk8<r8+S]���4،�T���;��G�p�*ߕx�^�`�TĖg�2�5��3.���"0� �p'��o�˫���6���}����ft��ύg�G?���-��M��lflI�G�@w�a�pÄ�r�!��%�<�u�5L��EԳ�_�I�Q�i�6^�x��d�u)%�%��C7�Oݣc�A_a	��a|m�9�w4��.,����}���o"�>;-QK:H$sd$���O��h�-%�Q|$oT�U��>t�@� ��S��oϑm����k��#���?�߮,ZJ��M�����3��~6p��K��ڈ����|���!�5A�"b�;OhBy+��z�����~|ի���~���#�kĢ�8��[�TD���~?���t[�^V �ȼ���t���|���)��lQY�p��P�ŉgv-- ����ϊ����Q�� �'�
��Q.���DKuX���y
��i%�"�]�#�d�*���Jk�^?����=@�d%LiC⯚q�L%K�<��-X�� ʚI�?�꓉��� �N��f)��WO���BtO^J5ff�@�����yI~�C�QfK�0?���"J�����}���C�ZV�P;J��ˆC@�p�?��9}2"K�6�m�n7�Oj�)6����e%}��|���@�eO�4?g�k�zk(�$�U�E�T&� ��҆8�cTH_)�K5�ōﺺ�=�E�����[��(��X"�\q�a‼����ڜ��d���5�w��^9�yy\QM�f��
�~b܃hI=п0m��ء��bοP�DY��a/�]/=M�O QQVB h3�H��fWŋ��b��3�<t�[�O̝�"H\lE�ou�U2t�{�V{4:��~��g�-+�$�wd�|k���`�q&�
Ǹ
�E�yq�8R:f�ԵYT���M���1��Š��H��mSO�9��i���'�moɲ���ő�����6����6�B����7������ԃV�;�Hij���K�PPS�q�Rqg%Z�a�)�|\�ַ��d��J��xr"���p;[(
-g�����:�m�]&� �1	�� �E����QQ[3���l��xJ_Hp��CA�5��!����t��%���/9���c���@k�A��/�ձ�/꯵=J�E5F��х�L����DC@��g��5UI,�9g�v �O^&��;	�&7D�����6�E�.��#��E�;�#^�\']���u�jce�d�94]�G��?m�e����^l���g��;�0w/~:nK���<�6mۯ}"0�'X��괧I�4��f�Ϣ\v����ҟ���,̋0�� \FP�,�j������o�hD��1��&�ۦI�Z��O�^�r��` �2��-�a0b��1�@��x֖vG�B��.�9�JT�&+H~��U8�$|f*^�"&{O�����Y>�q�I?�c2Bo?�;0ܺw?K�Ν��Jm�ܑ�T�w1K��G���ip�>�{9��,N9��?��u!�F�k!�b��)���3[�z�x4��h\���z�e�W��c��'��^�MMI[��I��Ǆ�U=��CU���E��1�GS�o�sN�����,�� ��	���f��'t]�.p/^,�v�o��?�uP`���w��E����}O����d���!ѶH�%Z�, s���&���y���'xTt�7h��8E]w7�4 ��D��3�Lɋ��<��M+�zWw��L��M� ;�YO� >wCϯ"Rn�aŇ�0EQn���B��#<�tA���\u�N�!��7ze�j���2��ё�U�P';�q�扗�E/��*VHjW�28�!v#�*b�����(���]$/`�´e�.������R��t8o�a�Q����g�g��j��65��J��t0<ǂAG/@�R'�'�!��5���@�NL����g�h�VgU�v�sō�ƈ�ش��OZ=�n%�T��&[�.�()+�}��MZ���8ط��a��O&�U ��|����҅�B1�9G�G�N��>�]�r����\�cۭ�(|�m��e�k�F$j�uϪg"�u�L���\���v2%�R���v}����*=;����!%ٝ!�����Iw�N�vi�ek������5}F�B�����Qz��N9[ژ�S;@�����6t#B��@o�C����ۊ��ݩcnV����_ϣy]�N!#�L��#�1�*R�?�ѷ��	l��oK�8BF	,Qi�H&G�)צ]�z/6�Q�I9`شeH���ӄ���+@�RӎT2�o6h�m��8�B�}j�yjߔ�X�}��.Co�#_E������g�*%��b�����Zp��l��g�wdV�{T��q��Q��B�X��?=� }�"�^��GDۡ�Ժ�"��rЂ��V���_��Gyk���r��*G�d$�~A��^?/����c��lK�(*c2k�aP�AlzBi�6v����g�e��\�(�w�.]s�r��c?��F~����3Hz��-�Ŀ �_z�}(�%�m6�Hx�lEX_��"��������!9�a��C�S5����+Z '*"L����Ә�c� fB�~�2���vn-w��S��.��ˈ�l��kyQ� �$�M��	o��/�:��<#�+Y����iؙ�a8�HϺ�\0B���W�S�Y��ݜƮ�g	fCo9��U��Y�*C1qG���y�J3��e����3<��i ����wǁ!o�Ӯ���rq����@�������T�z �*��ZXAVP�MӤn[x$\z�럊Sc��	�@��rµ��֘�%*h����j��8��(�<ҿ`�9DZ�H�JZWfG���1�r^�����|���ơy����)]C/��p�Llݷ��z���6C�÷�N�&0��d
͜�$�;E��{��B	>PCw���*>M0��'�[�͛9E��Y�dL�6L�jx�����:���#^c� gH�$�����E#�#x��x�R�y����0tU��y����#B�p���+��_q\��I�,vP�1�O&��DMO����l�n��)(�C�r=�8��><��,�F�{��?)HA6.��n�21kYX��T@7�$^qF�����@��Te)Ӏ�jiV�2�L�bH�I?ܵ>�E�	�-xG�<;6W�$(�<ͬ
8V^�]p�?��38?����+.=9�XQ����G���W�����%�b�D;h#I#�@��f[�cOp�3���8�F�v�c�Bu�I�#��$Z�c�w �p�>hh�w�4��ڧ`��!?�����S^ 2�iIv��l�P���o{S�^j�*�TSc6�$"���a���\��1�b4�/�]4b�)���}���5�~�y�
�S�cb=ѥXm�M��x��7��	.���1���4WW�j�����1t�h��?�":�#Խ���L OQ�O>�d�r��h�$�����?�Q�6�4����PW�$
��uN}��3������huX�rca�ݝ�dƌJ�w�D)k��<?���J/����w'"���w F�|Nz���=O��y] ��iWqu���o_ތ�<^��&����@�
�ox���>cp_�o˰���R"�8��N�����S\.��׍D�	8�R���hw8�Z�%t��j�ޱ�Pw{d�$N�C2�Q��Tc�t�wG����br0��~�A�l�l��.Ip�dF:k�򳽙:������P9"�PqlDǦ����3�&�/�c2+z�q�[P$��ml�]<c��|���ֺ+� ���B����.��	 �"��)g��P�g.{�y��.H��X� ���W��s���l&au�������9���U��p�M�3��2W�(�*R�*�sZ��P�`���^h�H��ߠP�w��%������PV7����+�V�P�l}�m�%���!�&vH���Pq�]�*[?��>��$��*��t�]X���JX�s~%[�?Kc����9��.*����R,�	����r�]3aVz��^��#�����K�tH]��(�#�O�����*�����HmXZ`�[	�4W0�]�`�%'�*��qGwGt����ĥP�ޖ�Pq��d�[��ږ�i���$W�[�vЁ����6&���7^�H�'�����ی�#,�x`��1��E�jȢMS�oJX�1J�#�k:8�W�C�n�[)�xȞh�n�ӧrVY�s�g1䓫�N��t�]�I�6�����K�qB��_�l,Rw7��D%-�l��m�B@�ݟ�yQ�~ k�_`�Qg���$�m��M!?{�ݕ��Z�Od��%�f<����?\�^��['1^c�k;(��
eɌ�C+jb�w���;
y����k����e(�4����w�.����j���
�jt��%oP��'��S�Wi�8�m�䨨�Y�?�pdv�`�~�W.\��3��Hk	t:	d�d=C��c��E����Ql2�����`���n��ؙ���|�6�/�X/�B�A�O©�^��
ˍA��bb�=��g:�z�jPB�3nG�Sú��e�;X�x�^	{Z��	��չ�:"��6������}ɗ۝���&Ƽ�B( ��}_D�b��Ft������'��x\��|)N�*�l�T�׃�\&܎Z4�Z� T�-��˒�����
<B�_2��"��
���dN�� ��b�j��'�u��}S�C�aH��gL&ﯱ�sVQJP�nk� 	��8�8�T��Q��8	g�M/�!$��J<rM��'U�'*y�8@ۨ�S?"�&��v �YZ��씪��8�_��%H����K%�
-N��\<!Lr�PU2�N�ĦF�`�кm�i���Y�]����Wq��#U!��)��E��N��SYo�?iV����k�<�tP���Ӏ�?�\A�¼�4�=�>6�����+�Mi�|}Ϥ��T�2;Mp���� �4��<�1x�2�`�.%�`xD�mM����C9��暫qO�W>r�PI�n1�0Ha�Z��#2���ocn�C�R��{���%�acN!�f�Fl�Md��=��`*�l���8�/��.�B��6�e�^�k(x���X˒��>ԯ����cԦ�y�T�*�ǥ���7ܣ oV5Fկ.c�N%��*�w�Z��
�c��M13��>׸����-&e��qsX��35�=:V(��F !�� �f2� 5�nNTMɓ���\D$�*~��6�؋R�:�t{�l��r��W�Y�Ns�%�?����|��!�>�6��C�v� ����� ni��XQ���.h�����G�}N��@���(�	�K��m��M5��۪lu$�wK����b���#���c��5r�{C	�~B)�C����x1ֶo��p�9�.��Ӎ;�Gs8#��)-����!��u&����5��Y[r�G*�,-]KMi��ӻ�9��7�aFG!��էCk��F�o:l\׊�0�9	!���ld�K����ç�f�,**m�g`v禚&Mr&k��q�8O���`X�
����M}��1��ZT�R����8A���)s�^�ϓ�������������(�m��P���Sw`ɚ�Bϻ_����������5����vtiڍ�� ��c�$��M����.`ԝ�,����t��ԵA����x^���8���3��;Bc4��t�En�6�R�u��pnS�3co�\���IC��o �쮮)����@�s@���u{f(<'9x2dm��>4���_���{�v�Ok{q����io%��3�<6���S7�D��,�fDtT6w���~��)O�Z�ׅ;ntPf�_�"!l�2�I/��r� ��V�  {�T��'�oʥ��= '��sر�}Sr~�����-Y�����YÚ{^����J�ꈢ���%����[���I��u�?nz@6�+�q�e�KQ*)8%ܚ�����̋�� �J��vŢ�Q)`��֭��~wf����+��Y�^�X��Qߘ���VFb)N��Y�sQRڏLɢ��!\��t�n�L�C�������N­E�>�H}}�C�⦙>{�!��.p�m�)ݹ'~���)���L��~�W����Cp|ãF�ۇ�5�S%���!v[�63x�	do�F:��mԨR�s[��T{,}>�ty��pq�0�z�l�*m�۔�z�1�W�� �KջV0�Y+։8��hA3b�ax���q�z�A|B��l�Eՙǣ]N6<������$��r���ER�65n���bJ�G��c��6H4<�P۞���@z���`��50���JvA�GOP�uZ���g�X�v�GoQvV;6�\?������yM�	4b�0%��t��W������1��C	�5WJ�U�tdهg#��
��
&Ҫ�pq蔺l�W�� �Kև�R��	E"o�����Y�������#�+��b)h����P4ón��i�	Dv�5ǟ'Pk��H�
��{n��u�0��Al�z�Mz��)t�L#�fm���`�l:Ҽ8�h�cH���' s���	2fe@_ྒྷ�Ν��q�U�n�iQ<Ӳ=6#U^�5�Wظq�1P�i�"e���AL�2�h�5𴜰���RZd�(�p��k`�ZBQm�F"�C����(R�����&���H��A�k��ńt��摯�m��i"��п���`i�����Kb�o�g�x5�3N^KoA�T6��q@���npH�^@/Ӛg	x<m�D1�������S3t�{�,��,��3db�-��a��x��&n���/ �`����Ez$����x.���#T�ɶ�������u�PW�>����?ZL�ɒќ/�v��ss�S]���c�4�ɿ������_�$�/�3mm8�ʄ�ɔS����]nw���ds4�Jఠ�� K�A���Q[ ~�V u,����.��MსFm�Pw8���`P�+�#�o�oF��Q䨎�̨�<��pkv��&V���ſ~ªt�h��P.1|Q,s.-*��ם[����*B^%��Eg`���c�(�L׃j��;�تV�by:��i��g�?�&TOג����+�*�Bo$}/b�2�d��
,���iN�:@hQ��Զ��GjQ��K��x��3���Tk��R���o��yO��i9:�Hs�[*Ҕ�XL�'��eɘƣ(Or*���=��:y��]�Ɣ�?[�%��z�/THS�8��F�ŏɫK����Ϳ$�F� ���Wns^A�?C&Y�">v�./�P󃾠����e߫�\�ɋ9�bJ�Gp����7�@�M���@ը�2=vVo�!��q�L���N�^h%[Ҭ�
����џy'���RMB����D�U��: ��	*1Aᴌ�\ �de��?��Y|��2i���.X��w�k��#�E~梬�_�@~g2i�A�V[���B�53�����W$��$ء^0���їlF3;�1E�O�].FPi�=�"xYť�E��}y��I+
fc'�%�Q��V���)���V��7���w�l�Y�����5�UO�ۍ��� ,�ނ����	�by}~�ݏ��K�˂�X5�)b�����"����Z�"B�TԹ���
.�эv�*��r滇(jh�i�y}���Jp�����@�'珲;վta������j�԰���(��H��Z��>�g�������j���F��R���l�ZW}(�۪)r<r�Aa/V��N.}g��k���5����:��wy�$����^E~�H���� ���嚷��t3�[�)���yȌL/��r�>)�H�j�7����^X��E rh�޴lx��Xʨ���$w;�.A�n`j]�y�Y�b�W�г.��w���!^�d`	p�N�o�����~�`Pj���s�-vxe����֊F���uN~��|��"v��N���/i|�.��b]P	�{���/c"�p��bKu�w�A�3@q�)F�7l��E���-��(l/L�j)CA=�v�bP�D��o�̠W���1���)�b[b,警�nY�á&呲�)8o�鲶�J�m��7p�����f�r;�Y;�u�~��5Z{>'���Eo�M��_v Z��dU1����B P/1xc����_2�J��oP�F+�]�������^	��ԣ���Đ��}o���>4a�S
OW�i>�u��)N2{[룇�	5PtR"�����\������x��`e�á�<I ���7����ƀ< �hM�3"d	,o7٫e�0�n��ίl~�RM���kBd����g$�e�g�GN����m������	O� ��J7����ϧ���t����pDa���&�Jܚ�������.$�&'�7j��9��?��m�����<����c����Ze̠~i�.��'���愖���,����;����e�՞�k�N9�
���-6ւy%h�͔�cB���V!�wȟg�QP�#~Jv�?�E��Θ/�{5m�^�PX��i��Oԏf�����d���H#ʁ�^��U�S�iM�� 75���C4-ֲB3������2z�
���֠�4K�n���_�ө��(�����}�-+�9��y@�C�(�A�'$e���p��X]�h�����옧��`V�fK�*�����|������yX��y9y�8�u�Z���V_��,w�J쨗>�/�����n����\3d�O�NX�YH��rvy=�԰X��^�o4��ˢ�SJu�0�p����ԕ��^R�?H����[���n"`<r��T\��XD������;Ԡ�����'Q�E�[MPi#�HMo����V��20:*k�J\m���H��]h������;3��؉�첓�œv�i�$�u��Š��^�&B/�@��ͻ���F�7��AU�e���}�9�� ��L�%j�(m�e���f�����]į)���(\�S>L�����J�4�:R]Aɶ&Yv&u�Cr�|�H��t`�����ͯ���1WC+N�{�����v�JTG(F7oY�ZO����ѝ��<��ta���o�$��
��Q�:�׽F�)bX����Y����x��e��&W9�V����H��r, 
��i��
Q�&|V����h1�E��Z 1�e马J0�(+M�%Z��3�J#�Y�p����y��i�Q���Z����0iV%=?`��ްtIP*��ljn�`;�`ɬ��dHn\:�S��G�w��-Wƪ'�A�˄9�%A�驡Q fG�>���-F��
�/�נ����y��|�hHn���@��e#����@J� �e�X�,�.��kqR�\M|�q��,��F�B�Rd�1�J��[��!�"[��n����Ƴm��3�v��%L�R�ӏv�S����� �s԰�m��a�i��_])���S=�ȓrY�H��nV��j�Ӿ�=BIf��~0@(�,�2�H�27�$���*�p�p�'^��-��O�X�HS���[nE����M�f��L��H�3�L����\�$a���2	e^.,��Y5冂�#���3���-��{69Rke"֚�����r��#�;F��9#^�L��oR�r^�Ԅk�����~a�I��5'G�D��X<� l��1���!'ˡ��&W1�����ͭ+�����t>�c�o�Ϻ�4�WC�"8��u������&{Bt7:ļ7uS�E��pʟ�pc3c��</�H��	�:Uз��1P�t�q^2�%,x���1̢�N����Ƭ�4d�&Af&�@UN���n�������*K/P�l�־�G�f��P5nSe���PQ���ܢ!��xJ��x?yh�И��H{ņ��UE�@Q t�Yfi���$��
(�
b2�[���=��o�E��{f�C�sH��?��?J�|����B��T�7��it���Qe�ꣵz��e��&���P\�.웬�1�N7K,�;�%N"G�~��@B25;u䦊e��P� �����j�rr�.7������l�|2�UV���!$�L��(����i�I���N1��Ϡ�,�����h�������5O*H�dJYmI}���[q�%С�S(<ux���	�c�tE?Ъ�S����𥣬�dApC�rn��vI�M�b��말��4?K� �~ZM{iD@���}���O
GEn��u~���?M��O�_��r�f��!���5����]{���x{_Ö���l��;�ۀ~���W�9K�VSs�ŖXkTC�		&w��UO!�v�
�,䰁��k|y�ɕH%A]��g�����Se�� $!�)��O�8Է��C�|�DR��=pf�]GҌL���vi~�T=*�4b1f�B3��%���<ˬ���f��1d?tF��:&v$�E�K"��t΁���Q�����h�	-�W4���e�xvd[�Cg��*������IBݹ�W�!�T�0��V%
�:P*��42lۣ9m;+3� �>l�Ut��Xt���ˬ�8}�\[es����;s�X��Z��'&�,���oE�0ij��=�N��ց��*0��CD�������i�F"j=�2_X����jsu�F��DS��;9��ѺT�+k��F��:�2h��Ip�(A�CB���/���Vh�T�;yw&��[�,��4D$����\Վl�<�)/����W���p�2��З��KQ��Ǯn��PywӲQ�R8�J5sz���6ԁfCĖ�5�A2_;.��A���
=eO�tz�1$?5��e�-ڃ	�� {z�ҹ[욙=�y�W�9�`�d򔗵���g׭6���L6V�S%���[�8}��(K�|�2��)wBtC>��_��Tا��5�w�Eǎ��T2T�Lݯ#X�rb9��֏�J�/%Af��6�{��0�m7 ����|B����.mY�V��v{n]��Ua2�Ö.i�R��9+3�5.E��5+Ҵk�sd�{vr��G��^�J����EP��I��YM]�[�&oAx����F��욲�+���������� ��4h ��hT��N�n�Җm��]��tAO�<�:��/o�����]$5}�Й��m�Ġ�U�%G���[*�PW���A�}�8���9���@[�*N�-��Z9�2�9��U��FA�l<#�ZL c�A�E6Vv�ǷU'T�6���?dk5��1
�Z$t��o���A+N��;0ݎ�E%��1V6v���ɑ[����O�����=x΍�G�?`�5�0lg]�&>IX'���l��:J ���~�cK����o�AH(6�%p{4��I#%��K�X�D���!Hy��#�8�a�OLk�*�;�DU�7#f��& �%�Ƅ��Gi�@�s�J����R7`O��c�,��2f�<<f����w�6`ޠ����MƯ#|t�߳����i�}8�#X��?Sa����H�5ش�qq���j����V�_�r��^�eo�C�9!�5	��bnު`�7�I::	�66��f���0#x+a�qLp
��nD��+(���Py�We2�LcqU���h+�feNc��ĭ8���a�Q_rPej�VTɠ�E���k�����!F��vL�i��L����[l�3���@�������	3ǦUf�ɤY�-u������&��׮�o%��S)_e'���a�=�_�t���y�@Ќ;Z�,�-��l�_��QD��B2��/'\�-��mt�f�O��ը֓�DU^F+EzFK5�Ϥd���&�m����/rm`IjvKz�y=&��h�%J{+����Dj�+�A�M>O�6r^$������on��H�c�H��ޢ���'��v�q�Il�Oϒ�]���HK�F�t<�XǬ�f�<�5��-*��Q��\��ce3k�H���)<�S�,�9���5�?)A�E��5{���\r/v�/[bo�LE��?{��dş=��[��\�x�H��5��b��H~g\���&�N�A�{��!�o*��Ne�AO,���Q1�y�F��S�i�O��u�|��7A����Q���T�i,ƈ��:k��a���)�.[����S��ɒ��44�e�S^X�[/��?�X4�S�nU"�/�:yPI��]�ў�oȔ�5Κ ^Z��u�핟t����n�_��Ő����v��Կ�ɇ�"N�K.�4��<��(���&edl��}��㱻����*h�䥇l��V��<2n_�ԅ��h�>���BC�&���e��j�\�ݟN�>�HU�f)x�G���f���z��N)���}J�6{��`ҟT��v����v����o��z����!�7�_>e�P�ф��qG�xTR�k���j�W�H�ߊ��p28 ���+��W<���)�Gܐ��j;0����!�(�+�K�Z�B�M q��뎲\�qm0^��I��~#4b��=���Jʶo�d�rPOD5��rp���Y^,�E�㧓���0 `uR��:�
���ԄF���]����bؾ��ۨ�l_��/��R��V���V�(��aTGB��,>����p�� (�Ѿ��w��O49Ujh�,q�xfF����W����%ǐ�dH7şeE�5+zK�Ț�
����<7H���@Ԏ�F���������iȘ�յ���s1,������?|�Szܻ��=�RR�e��UD�X��c�9�]�
k�:CSa(Uv���d��Y�b��[�[��s�A�C���c��a�J��c��]�$L������B�����WX"� �qt�4h{��e:�����؇g� �c��g�gy>?%��>U��V^5c�Ah=h>�� ��[�(�w���Lv�|{���:�����n�lF�zj��S��� Q�����jg�t�3`��h  4l�S{P�R���E�`���%�!S� ��}���h@��3���	�3�S�ej�e�lL����_�E��v�[ڜQSuDL�K��xT���e��X ^��7��s�U4��O*���T�����̾�� �$�G�CRt5�8�s�Vk���2�����LD�3?V�q+�U���X�h�j�u��t���Y���'']nm��׭Y��v�i�_XP��_d�H��lXA�$�yM:h1��>�(���lt���,��u��}8��n�ƍ堪TCf�:~��|㶼��Օ��^3m��¯��ȋ��q_M� ����/�r�E*�+�?��LUn����̦��j�����nsp��<q��氍vkuĬ���pk�֙@�L+���s(�I��S�8p�����^�#�dU�S��v��b�z�s_>%L�L�&��ÍW>��[G��m�HO����`E5���'�J����8��Cݛ��E��j�ǹ�>}�W��A[�'��#|��)g"��Q�%R��}�j���Y,7ѺF�DNi����īm���B��,�x����4c�~�ZG~HX47V�l�3l��xjo\Q�����B�P��DV���@Jˣ�S��ϴK�^�̖@�N��,Lt�����3z�_@����<�����Jx�[�wm�������bRb�J/WwbP�����<��l��|,䧗��(� bd���i<߹?�eZV:�D��n�U�84��䥡g�nr	h�d�	�m��'IZ��b�����2�6�O�8���� �Rp�gnP+�3��rZ�
����.��y��!<H���O��ˈa���i8R汵#eT��>�4����7�*����4�����Ǡ����Y;�c������awS��AѮ��g�l�r�-p�^��Ϸ|*L��ho��Ơ4���-�#I�D��ox&��,
��-���D/da*ʅ��A)��n�kf�CO^��f����FbF��f����x(FAk���[27[T��=W�g�uX��&� s��1~"�\��?�}瓉�p�k�S��������k��{}�L.�vP-raM�QLmw���F�V��r�J���:w$�J��<Y���R}��'��/�L:
�a����Ng���m]�6H�5�V@�uyE���j	kms�����	92�q��GBՇ��
�k�d3��:>cF������d`a�nb������,����]�!�1��L�o��,�\'��/��:g��K탐�[�����>�C4�Yxľ�ԟ��Bv#U�> �$�nRg!��� �
C�ȧ}�Ĩț�1hq\�xY��JS��n������h����}Y�`�iih0]�(�
��4�E�˺���.R��M�څJK39!L�7Kw��� 	��ۮ%&��ˎ��t���qn1/f"��\*�^c����{�m�)#�Wƌ_�}���si83��^���樣�S3�Vƞ#�� ä�7��<�XKI#u>;���h�%$Ao;r�#��.��0�a}��BV�{�]ĸ���O(�yny��������	l��,[�&�92e(�\[��v�w-�!�&�}yj>f����i���p�"+� _��N�vQy<rM�	��(�!�Fm�>���w��D<G�ǁ��8��e�&M��Э��ˇ�L.5���v]�ؔ���.��}5l^}�"e��)̒?�ǥƴ��z1�����ę�u�)4�mC�_"��3o>ٓ��q�~t�^	�����%��l:e#��z��j��6��p���;:�Юc�.�O�������HU[�˺(0Z1"��k�+�T)2�G�!z�hm4p��87�0�D�dX��C#Ǫк���rf�qs����'L�~�L�b3Ψ��/��=adc��q{&N���r���6)u�zG��{��^�R.1���+s[e�+��6t ҕ'���J���t��"���9d�?뫭x�h��b�(H��<�Y�4��&R��W�0 �B"�+n2�SZ�4��$/���`ފ���j�cu��m���+���e����pb$�)�U	\���bp)�Q�j��znS����á�9`����u��Т2��:���*�\sI%K����7;�쀤��;z��7̦�� ���K�jc�wcsI��/=4�6������V"u@��h��$G\(�[�NA"�Hc8$�\/B��T�4 4ck��\�t�*`\�����L�7�Je�/m E.�Z�d<))d}�VW�� �3�t<����i��}��M`�pI�F�l����1w�וNV�-�(��_k���{(�~$y�2��䳔5Օ�V<���Q'U@��1�9pK	Һ	<��q|�I�>�5��Α�o+#�Ú�C���(����Ró5�
����M˂u5�'���u)�W��a:.Y�@m��r�;$�	ҡ'K��P~�F��-:�z_k_��Lޠ��� �i^p!�S&Pa^��r`M�Yn�*-u���rU�y������G�S��B+�y�*�9�ٮ��d���,��8�֙,���:f��Z�Z��U�g�F��T-��x�Á�u҇�.)'������As���C5ik|���4'¦Z�����2\��ѯ�}�%S(SEכ�h/�{�K�w�K@u������Y��RJ�θ���s��)8rY�6V��ԼH�o�=�8D���~�����@{ə�Y͙ؓCd)�>:�w}��ܲ�f]Pe;+��-O��*��2�F�AK��4�$֘y0 QLqm�Dp;�Ĵ��n��j|R�ߒ�]Sw~R��E�M@�-�-J�S�L1����Ad�zXyӧo��N��­��[�k�Do:k�,6@�q[����}(9�r�YwUFC�D�~�Ӟ�!;z�:��n�DQ�P%̩�/,[w��6��KEa�u��Ve�!0��'�DB��:�$��+�����ށT®��X�M�oL�ic=�On���CT���]�$�r�*��B�Q�%�������������D�G���Y����_n�P�  �f��r���u�倏�:�\K��� �f��ր-�a�?����phW�m����d��3�<>�� ֬!�n�o�	,�A9:�y>���`�3�S����v��/��IWR�5�i��ȶ��:����0۞�{��7`����kV���g�I%��Z{�ẅ́�F��6�L���pz_�/�hzm��{�����xw��)�I|��ﭹBIH�x=�'�ٺ�h~,����)G�K@%j��|y/��T�3��_F�ę�|�ƈ蜶&���"�PC~�f��Vkd#�`�$�4�v�z�X��׉:��yGjh"�eO"v��&��R�����5>4&��^�ޱ7����j�8q�FI�_�4q(Б/��O`���ґa�Z+6�Is��+���V ��p����}��ty?k�`]0���h����#A�l�5S�?���JA������DJ��g�3O�@᣶�B�/VT�tZ���>Ҭ9(T����0��+��{a?�Ύ@��Ǿ���7�_݊���z�-hF����F�0^m!�q�X�fIng��^)�Ѵ��#Pݧ�Qv#a7�����p��4���',a���>v�x�c������!_��K��6vo���-(�(�f���h���p	<���������`�_ ��(أs@��{o&�]1<���6�/�[��cn='�bo�5mH��i߫��,����V,�p;���WХR�`�p|hoi��!Pڏi�`�2��P	Ϟ>~��B� 7�7���(�e��!�q`�R��{ȃam22�P��G����@�!Y|����ߚ<k;�Jd��S�,hS�n���0?��k+����s��ߑP���t�H�{sݡS뗞0��ْc����RE�h`;���A��aI��M�I���KJ�W��C�(�T�ϡgEy��I^�<O{r�0ՠ__�׷x��0��6��[b���Qt��$Ke1�9@*\��i��+~ܸ�P��CJ�z��}�������Cĥ�
�BB8��^Mw�S�C ?'g'��Eιt��;J�������ol��Uwج �e��7�A��?^
\��:Iҽ�/%�(A/M�k�#�Ҽ�g�Hv��][�.ffS�Ka�%+iɲ�?ta$����V�(N��	?�C�z�L}l�v��\��W�����@�Ch]B��×BAX�+ 3�`я2��%�8�����W�NSE�"����(s���I�M-s��f�ǃ/�s��N�C��q�D2+�t���N�^
޵���Dx�}s�M)�[�u��6)8g��r�Mx�Q�ː
�$��$?Y�?_�,�cX��FR�����4�H�{@Ȉ8/�t�g�BwLE1�$l��X4�*9м�%�ґ8��ͮ��A��G9�4��O��I,��=�{�1�\6�$|�:��l�a���~fsw[#��D�bN�ֽ]M3&�WӤ;���픶����v�kG���`��y���@G�#ٟ���Vyu�'nc���͇�<H�(�8o��o�����.4	YV;�A�Wr̚�`���C�e� u	�%]ÎG,�(X����������$�U���W9X��t����.�`�f�2I��celu�-�e��Z�t4����ުk�]�Ι��z)�_�j���������t_����C8Vb@H��L�4m��� �Cۛ��`!�:� G�?\�SO�׍{���� ��W��e8zj��m>]7T�,��x;9�}v]v�0ץŷ��k2���XFwa,?q/)�YC�d��'2���Q�q�<���`�kG7��.7��iWKs4(-t%�'�,��Y��7��%�I����>J���e����G����S*>�s�ђGY)CT߳�s�h��OB������\rtC7�=i1�Kr��vWL����	21����p��DZ���Q�v��g�J2؋}��ӹ���j�w�w=�~}��t���q����y����#p΁��xo��ގ����YŴ:2�꟏�ڊ����T_�s���/�@��z
juep~��{�:�V�0M��t
�8�6�~ybY�P�>e�X�,/�&E�A��N�Q�C���B���[a���B!~��$;Y�b�\������~�p?�8�0�4�e�2�7��U��Y�Z�QS��p�������
��A�W�~�״�@�4���q	u'@��Ra��z��%�l˷�Y�zq�lʽ��ƴ�L�^V\�?[$H�sx`SKi����|{.M>O���_��r��:VֆဏBox`�Ŭ@�l�%^����r�B1k��Olٿ��Q=�"�T���ʨL����z3�u��:��@���IP��V���@�)�4q��F��ɤ��5$���7)a�w �5�����N�B����bg�����L��6��h.��j n4}9���:�<����TyH�3�Q+f+��,HyR���ח�a(O�{)	q���f�7v��0R���O0�EFQ��oHu����[YQ��mOf{�����z�	�nT&)�M��YBE֗X
�|��M�@�.��E�G89h��q�&oX'z��j�5�Kr�rQ���:)n�_�H#�q�kCT\7'u��Ϭ�ò-�R��`���[�d,;�uT��/V�q(=�'���j��VK�e��oHd��ɵ����.	u5I��%S[��#v7x���%�OxDY�4�m����#�ZD �ݠ�$5Cņt$R�KkK�r��U�/���Z�[`��W| L������ǘ�b��w�<�g�O�!Z
�o׾'K)�9 �W�1����fTIe��J�$Ϥ��oG�Q�SS��+F���+�HY�U��uG�7���\9~�$t�X�O�g�8�Ȫ�E2�b��s��]%���I>��pN��R_ n���7&i�ނ̰�~�J�O����Cc�E<7�I7E��Z��뽊\�I�*;�����z�jb��zK���r�]-H�>+s�xtC!3��S,1/��F�I}|�(��ٹl͠��`��iQ�c�,�)��?��N�־��Y�n4Y�˼d�ls�h�|6�/GoP�=t�<��Q`��im�%t-���-���vu�J'��;7��N�Y��Y` �����H���}���k$'y�p\����5C?I�L��o3�(!IL�Ej&e���7�q[�F����fH9qɼg�/(�}����nӍOjT�EJso�=�y/<�{]�z��9�[4!.F��D0�u�0������nb&�&5o`��8��U�%�8��B�?|���yt_�y�Ӿ�J:���攽�پ i �7�� �#������=~�֧L��7p)��	"��TfN͔,��r���7�1���@>;���(�	A��"�+��gm8�m.��-oy��K(�?Q7Ѝ,,.w��A �=��e�b��x��s*;.J�|�,��4aѹ������`�=7���
EY���S�ŮO������Sӣs��|/���{<�ʥq��R��:�V�:ń7��3	�t����P���Bvumb�V��4�{j�k��k:�N���)kԜQ:_��㞂m.����&�����)�/#�E�#lo�������G�aK�;�̰?��e��W
�V�v���i��l�� �k����Q����6�����>���NtI9�����,�ޭ�Z����|��q��*�y���d���:6�[�-#�+Z^�:�~�M@q��HŔkh���^&��X�@�nN�����1��O�P��i����uBML�N/�E�t���W��G����_���r��o��cY�o�!α�C?�3곘�]SyV�)��O!��#[w)������V�=kb�c&�J]D�"�Ɖ�N��di���NZ��_�Am��ge�C=j �$z�|&d+<# �!�5�f�� ���1�CT$/�r��k�cjRd�^��y`7��M��۽̨/q!�G,bGﾝn��U+���0��7k}K���G J�ؚ�vHǨi5��ɚ�=�7�JY}=;���ed�c�-l�@&q�B�g�M����C�G>����qτacQ�7��<:���n-��'�[��
�RV.�#K�U���2|}֡�5�J�T�B�:�r-B֛f��$
:�ᖂT� �Y-hY�d��Rc�V�*���R��g+!\jLB�Qn%���IūW����Fq�?��X��,!�y�t^	��s��q�,e�@�f>^}}.N�b�Az�7�v��Z���C�W� ]U1j��Z��\h��̭f��'Z|��r�0��$�����ҵ��?�ڴ���I��c�KW(�P^mgܤ�W=�� �Z;���{����ދ�љ�-XtYLgM���h{5�	��}[qݘ蕮����]��7o2��f�i��Z��Y��i���.��w���-^56��-#�_[�s�F�y+���>SJ��E��s��� �31W�fܶ�����F�;t+[���CZl��;���(
�z
��T|�Y�.��K 
���~S��T"+zb�p���&]�@�f����Zm|��QxQ�*���0�a6�BT���Ԟ U&h]#u��M�m0	4�����+~r'E��Eo�x�?�o��ѐ�p�_�i]@��!Q,��y+8�+�z��B��4�����W y��7��^}��<�ģn�!�A�Wyr�x�@�N`��wY�3L�c>��������W�E���C͕/ͻ��@�qj�Zv0��OR{׆���01Y.�L�.��C�WOa�d��o%/A�K�d1�;[D�4��U��Ŧ�w��vWp�}`�k������̐ؗy��L#����ܧF���Nd1�tu0{�-DSL��k#F�tp���T�}����$�&'����n*|��3@3P������ԲWD��
�4���K��Ï�d���*��	�����k���ԘG�b�彷���@�	����Γ�j0�J9
$�`j��X��"5\�����d����C�/?������x/�3>j�f�`���nG_�g%���̦�]/���u�B�1�W|��h����M������j�%�!��7HHV��&�#{���_�O��-ǽG����2G7�k�����xR޵oï������\���G��$p���o)E�.�LԹ�kR�i�Szο0Jnsb$��Hz�R4�=����;S���g(7�<�g�bX
���Q?8����牎Z��]�|�&��a��pÜS�~$s$���"W�1gS��� �����R��i���i�ПD��c�~���|2%�Y�ٱ��ɽ�%�v��F� �&�D6|�ͅ	۶��#��w΋���i�2'1��闥�����Xx `w���s6Z�룒"��1��،Gx��ɾϚ�����KĢ���b	�f��O�L�R�ܕCa'�u	����D�e�u � g)�PW�q�.��8�[��U�e��¤ �Be�U�FQ�s�T��=��Š(�8�\�%��c��ƁXK!���6����+���a�� N��2�#�������:�]Ė73k#ʏ!U⦒ �6���+9��z+��^�8eẾ
�*<A�*GZtH:�ut����N����6����2v��?k��Ǜg�ܺ.㐔f��k(>e�lL|vm@y|�s��δ1���i��<u��{(������@��C�?���W���r!� ������E��6�z�5J�����8��f]����) �q��K�F
t��m@�e�f���h�ɶl�D��@*����d�N4W��b���V�$w�g�x�D�eJ���5�E�g�b.�4�[�0�����'�n��)1� P�COr�>"0w�,{;^zE5�̨���X:+?I��mn�[��Ӧn$ ��q ��Z�V�yjT&k�����Y��1��{��C˓sd�!	VX芁�s��<���R&�p?h
�������O�����&�[mP�k��w$φ�2����dcX��J#F����۝�vI�e�,	[�Z��=�)�Ly�ȝ����P8
|wE @%k!�J��"pD`?���+I�	*���&�4�g����6̬�����������J����ʽ���Y|��^�e�p]!���_d�f:Ɖ'u�)W����I�{)��;7�;k{*��\V�c�A�~���f=�O�ӑ�Rl4�<̠{|��&��鄚O��f�ٲo?<�����O���Ds��xCx����BJ������$Q/_��Z��/2z B��g�o�skoA�Z�lo����9k�$u\[�S�S8�M��4���p��]J	H/�gt,�����r�`��ʬ��~.��O��ME�w`�^��hW:�qR�o4u��-p~/	J_)<I��.�q�|4�'�)%�x�h�.1C����Av;�5v����LOW�NZE8�)=g���~]�v#�(��W+�c��M�6�$)+վ�OvQCr�2�[@ZN0� ��
�#t/�r��"s���@>$
<N�K� [�~��|<�E�6#>F���ug�&�Շ�*մCcVh��y?{C��Z���^~{�{{Ք��-�����KɸDכ%WE��=��X_���GD}�ږt��T=�0b��1E��a���ޮaX�'Qq(��н%�͇S�K�/��j�Vb�90؝��/��l-$��"i��\�ޠz�w�9���Q<TV�_�DI����]F��Ϝ#?���mԖ����9�hlC��uH	�!F�D8��4�}����IZh���)���C��hO(B=��{�[���O7���+y��	@�{Ǻ�؈�� zxS�L���R��}3��`��kkֽKn�M��6������|���4��69��[C4�"�-Q���<��F�}�N��5��"{V�g��rD������=������G�	ː�r���Y�a]���\)I�-y��E1���R�34-&_= �`�� ��~	�4��d�p�s������uK4��.����l�����n��zKf�v%j���iv�y����>�,=S.w�HO[PB;���5��ܽ����`J��������N�j�T�^��G$'�ZN�����q�RA�����Y=;{1�n �x�7�1؈u%�CŪ��XZޤ�(W��-i=��qkx��`kfb��7����T����r) L��k� �o����MvE_����,oԫ\"�$�^ �1���l���«<�ܽ	�!��Yy�<[�\�ԧ߇ڷ�1������	�����E	Y��2�v�Jm�a��ȓx�X�K��\��1ǟqv����������9& z�Id�}�H��Զv�G�:b��lIg��jW�mb8ag���k�H^[�c,�ٱ�Ʒu�h���C%(�{pZ��GO�*����cj�F�gN���,��Z���2����v��"7찄`^���9ؐ+w�H�U���w��V�6T�!���%i����8�3�ZJv"U�^���ੑ
��W�qr߅%�.C�4Rz�3<��7����Xla�_D�x��n��:���R��(�%YoW����_τM��*�\P ��OF\��3�|b	>%2V	��6�݌��<#ُ�zJ����,VF�ot
����7(���}��^�)� 89h��H��$pA!]�{���23���";��9�]����Z���u.oj����#����m�P6"Э���7�E�����9�s	�Ͽj��{�۔ �����>�!��đ���9�DE�Q���:�(�6J#��F%�p��x����5������R'	��;أ?�9�Q)��/��F�
͕���&k������� i�[�)P��H��[̓I��kw>1ɾ	�y}��WI�s,�N��E���E1�Yߟʖ	[A���'J�_�8`�|[F���6ɟ��f$G��u`�%�WN%�?�����ةC&5R9x[5�/é,��%H�p�gX6�	�����T���U�۟��.~aOAy�_��-�_~��"�U�+�p��qz�Φ��
.�;�<�O�t�PRL���cn��_V�[d	��e��wvM��KD3�)v3.��F��g������2A���uP��SŃ�D��Yˌw:3r7���sY�n�M$8�����IO�*�����x�G"�0�%|a�$�#F���)q���7{3|��F���=<�=y�v���0�F�����}=;F+#Bջ�N6�,E~��;l��L�� �HO���t>u�Y�t8X��	|��9�e���mtP8T�o0]g��{�#},��y ϥ�ږ]"b��c��R�z��Je) MQ#����\���[V���m_%"e`���	������(1���,��I=�!҅�R�aj��44���ZMF�����Sb�m�{�;{��L˱��1L�b/�M��3��.i.k&�����/��������cy�<���P}=D��㰖���k'��1*p-pHC��,�L��\�Mvz����f�Z�A�o��:�<�����p5!����؂J@�g��qe�4�OP���N�cJV�r�w'6�FN�fX��.�+Q�<���l�.h�tIp]�(�S��/ݧW�ϝ��c|�$&*����=h ]
��n:.颧�99\�I��6*��Bd�Z䍥���_ざ Z���[8޹=�z�#� F�\Ӟ��E�jb|�'��S1�9 1�2y�7)�N��?ռ$R���� �� r�g�P�M�h�ZO���Xo .#i�������QL)�h��#3�*�y~�d��<HQ����8}��dg���e
v��#��TL3�q��]|贏��.��I8D˸.s�](D:x�@Z���	�&8�cU��X�@>3s��Z�Iy�BH֌����o��,��;���K�M�d���\}�9�����U2^6���K��2�S�ˊ���q��=���F���v+�p�o�I/�P�gu���C �<��=��W�Z��f�=O�0������f���+��Z�����UD���ZH�s!Q��]��V[�ǯ���U���ى2�o��I䮍ʚQp̵9��.;�G��C]�Ɖ��W�A4(���R5�� �g��id�̧(�L_�P�	�:O5t�Y>u�^��.��y�,r�?�O����g�39��i9�uxw���lە�@��~:R�7�qh}�s�<ߩ�q�a	�A�[���R Xq=2�����G���njC���<��8�+ݙ�B�sW�95�Heqx`/�=��Xކ�=j���D�cA�^	���M���������և�a���p=}��ǀ2��W���_i���>|�x�鈷�Z����޿�|���|D���p��f�-�]|p�h�����fFÎP���K����;��Ҽ���<e�XKb��5l����<4��ȸC#��L�"�OJ���@��KA��P�V=ix͵C��l$���f��-W뺠؀a�B�ͼ
r	���~��+����|��L	_��BZ�0qt7M`�۔j����;PJ��
^�����J\`O�])y(m�X&2�(�H�ӛ���ox�X_�4�Sk�﹨f��M��I��1��7RNi�[oH�r����m F7g�>"j� BqD6E��
o�[��w��#�G�"Ŧ�ld]�&�����$�#Q� �f��,1�fҩ>J��2�G�'�����C+���^\����x���X>a�`�N�,���9�hʴ�H�^����e~�ڑ�����c�'!t֗ H��	,����U�_25chr�~u����Q��R��I苼�|@���?�6�gʴEnJ4���4C�';�6�E��1UNK��u�(��(��� ��6Г7�v��I���K����hі��˻�%��K�Q���\+>��6��Ж���yzp�Zw)-HD\"MK�A��:�b�н�R9|�rs��v��*qEy���}Y�:da��7\��Ħ����oĶW,3��zx�T�5 �,�cVnF�K^�b�<���u9K=]��?jQ�#9z������h�Zc���-�>Å����^��.{k��.�+�#��Þ66���]���s�;V�ab�=���˩���d�?CMM�Uݕx J%Wq�k o��-H!
,��)/�u{�P0C��N�CN�Qzi" GW�a-�u%鯖|\g�m��%
J���P�mu*MzK�H��?�Ɓ��x�6�Ju�4�1��F��S���r��o3۝����%Dd��q�ŗs��EZ�ǫ0���5OB�g����7��q�(KW6#���������Ʊ����8�CvMNs���@��!�Fe�7�z��#�8ԙf�t94�S�:M.�([[�~�w�~����/��D���s�H�y�bd>V�����{���|���7�8U~�k�r�����%�c��ye�1E�3�r������	(�
�O4�%�j&�Q�a��j�t� V�,����YD��slk����b��ή�o�|?�!������:7W��6]����m�?A'��.�(�C	A�}i2�u���P��00�nd|3�I��m�� G��yu�x��ƾ�b!���q��m��mo#��.A����I��D�������2����&:�%����[M�o�v�:1ݲW]���0mN�zjU�M(��!�=�֣���Qt_6�W��U?�1ՅF��y�׶� �'�jT����'�hC��k�A4���q������;�T0R�F�-w��Cm��Ǵ�X:��2�ˀ����C��,!}vu��y|;��v]��wv�Y�t��'ܑ�����d���n����-	��
��H4r���cL���R�ϯؓ�2� ZJ+���!&���v)�l��qZ4�&7J�==��L��E6�H�G���8����Qt���(�Õu��� �ӈ�$�ߏ��{w?�����������,!�XVֹ>�ªź̛v.��6 c�Hbd
��õqy3�A�fNqSz�lU�Ew��K�n��Mת�X��������1/	�y��U?�V��������Ti��,p�z��o(@�Y|���up<H��?LVW�!��rǍ��z3>�O�@���z�Zo.زv�W���ƁQ@��}� ��(��i���P��{ �h�p�c�DTd�.'5"�%��U�F���t7�լ����3�⭥_���}����m����P�������KzF�v0f�5�i �_��t��L�̔
_8���U`2�z�U��'��eޣ�[��V��[Ն�j�E�����/��n`V%��s�� ���n��^)���>)�)�����9���z~KP:^b���6��^�ܭ�*K�*Nx�H�Z��VT!EF�U�N~�d���x�[���j2G�c�q����]H��I�'�o���_�_���	ǋ5�~�\��%���Q��)H�s�f@���S��Ц�ri"��*�q�7W���L�>��j�����?br҃)>8@��iX6G�2���?5X>`���[>(�Z1�v#0�o�k�z���N��ظDS��v��|���s`>�ퟬ�'�����P��YZn�:��B7�6���^�Q�����a�/��$��_8��U{Ts�Q�k�rN���Yϐ�As�s��|�d����wV���,��`�3L�^�I�^��M�p�`���wSj`���/�ϭ^Md�4�!���ȅu��i�ڇ;�ǰ�ɳ+|x�m��@{�\�)�U�P��z��tk���P�+yّB)�6N7�G���Ac�<�%�1n�m
��J����.�Y��$0���h̢�����*ۉN��|��d�lVޯ�u)Ċ��:'O�4��c-%?�qCy������E�yV�����-�B�S
��
v��w���Εt+єu}�Vl��5���!��,�M��l7��	�
Gd�������������ߞ�s��L���P�F����%��������6��O{�E*��GV'�v/����'��X�%���H<ng�#��W� E��Ȥغng�|z/�.]~�:u�&�n��-��N���`ϓ���7K�E���hs레�4���n����rH���}]���9�������s^��bs�]��y����P���²W�g�]��A,�@|��� �N٩���C����#�ͧ���*����(�0�Ϳ��8aݽVi����"Y=}Z���M��� 6�����͈��ZS�_�H!![R�'3�ln̛�)��P��AJ\�CL�J���X_�se����%��L��hT�o�:Ug��	�I���4���,�����U?�i���P��zy�	�ᖤ�m*T��H��> 6Ֆ˿D�-��Is�=��	;|[��4 _S�-¤�� �2�����U�Ӷ�����1[VR/u�Wp7�-��� 3d'�1MJQ����<�Ɓ�[װ ���ۃ��d��N'���EC�����^��,���Rz�שf�����'3�vߕ�0�E����p>��=�0�6U6;��:'w?�v�����7P7\a�vt��]ZX\���$�$����*B�u�6�8}!@U���ܐT�Q���G6>�'��M,z)P����C��a'��]�آ4{?tOV�ǥ%[��υ�^�2W�^�ޒ� A^*c۾������Ը�ACA�m5V���S4[��ů=�w��`�C�#�k�_��>����w��Ko���F�3h���]��=l�"^�?�(�-��0��dArX�
�A֤��j��4�u�10a�.8�+���G]l����_w��)k���@�����l�p��B�w|��T�/��/������[�p���j"��A�)90\���y13�ٴS������IH�2�͟L��$�N�]Jl)6��G�(@Rx�9X	���Ɣ������{�U��T�4�Ƿلʉ�K����!3�tXai�E<��;~��(SOٚ�Ojo�>��s�����*)>k�ѸE�1���M��V�Y�)��0Kլ9c~��0������&1��m�s(�9����^ɦ`�G�J	���C[��4N�1|[y�&8�o�2B��u���s�\�z׃�$���Um@^l � �yjPw:F	u��10�ˌ�;�A7\P)�b�A�/i0�Z~��g���O�-�q�Q�MD��`��n�.�]5��|�5�P�y���ϵ��%��OV������"�-n]�+�P�!Z�����?�XM�V�#t��S�!�G��	0xS���Ҍ�U0�����~��Y�y+gW>h��!GBD��P��њ�2H��R�x8ƱR�4�'������4����m�d�!c�&_�I��� ��"0�d��oI���5��%?/����E�:2R�a�L�.R]Ax���b���J��R�nف�o�u�{�Q��!9������r�5`�z��2�%�H����e���gjc���7��y�))i�j]�x�{���:���"���TY.J]'4�²�ų�5� �W�GXn����#Izk�%���2�U=L
Fl��RO�?9��(<65ö�F�i�0����,-WN�X�tUD�n�˾U��*v��F�Z��RM��vs;{��༅^-]D�m4�ó�1� F��5|�m�̬�s�Cl{��������b�t������<�X�%Q�{-��ل�5�%.�sԗ"?[��������O=o�I.�l���Ԍ�������O���06<�<���A|�.��?6�
�[�+}>�W,qV� W�PU�q=i���b����:/D��D���د'�o�"��RX���ӊ�������Ĭ���Au�R{�Pp��Ó�����9���)�.��x�d�ƴ�|N,�I�QV�������s���ֆ�8��zx��]�������J�y�(�!�3k�Yi��CE@�+x�����������ޯ
ah���\Y�(d�I6QV�[��øM�݆�oc�m�P��_>>՗�.�2��j��
�����f�ئ(�:��[��J�6�^��Qp�	�W���������{u z/~_�wY c���z"Ta[�T[�0��4!Jo�oB�K��@y���Yq�53�hC��O�:ijv���Y~��ôJa��}|c,�Z�����9n�i����o<����]V��~*������~>�ɺ��k,/��� �7E�B�)��r��1��JgVO�4:�x4�����/����0�3�8�=b\��� S��h�$��iМ:��n��	7�G8��	�l��f��)IL��yp��Xk"�ka�OMi^0�"��m�z߼�B��)�*��D�9�M�;)���_�l���\.z�Yֈ��J���r&�~���t���մ�����!�9t��{&��)i��- s���\�h�T��dݚ@���q����d�[�Dv�2j�ޓ,Si;l��]��Yڲ^�����۱��+2VsB��H7\�é]�ޑ����j�Q��<HA
Gٚ��|���)�r� �µg��I���Z�3�I�<=�^v�=�Oc�M�O�]ȿ����-5��%;O�n��mx��i<hg&v�j`x�[�D�8��D����6��T����S����E�r��E�3��&�CJ���V͈��rvD^��V���E�R�AjU�(���یq�O��)�|z4��N�,U0 ��m��^2ϋ!��m}P�V��L{�h�d�~@��yw��s��5c�?�'��d��Z 
�0Z��*��2793TVf�df�ef cPib����T��cn�cE��,�\�����٣�^����_�Jβ{$+1��+qc5�;��ܩ�;�`b���ӟ�J#s�]������SmX�ڂ��2 �6�7h��x�8a@�LuC��U���4KX��?~�;NK܀��ۿ�'��� QV {�VQؽ���u�
�ߺ�gm��1v�j2�<?���aoc�Wye�(I�)Ҕ�6�w����ü���Zl��2�8��˭	j r�W�Ia�����YǙ֝��+�M��r��G��<Z.�zl��W�"1�RX�����:�m����
4�o/�<�l�o�u��]��$�,ߩh,O��N�u1EL�2���^	[+
��?��9xG�؂�L�i�+�� �_��`��nuz����K�ş��XgE�N��foK���	��ԝ��orΜ���� �}7�M{O�E��L'@ϊ�/{��E���L����o���a1����n��M^i�������ׂ`~������0�_T7��])o5�����s��n��٦)֠>��I�1�[%�p`{C�t�L!?}+?_\	��u7���7���.���a��4�ư�5���|b�Hv�[&�&�8��__xɏ�cZ��y��e�X_7� !����Dʱf՜�o%!��O���v5�r��j)�<9��<:n���J�v������i7�گ��+Z�����x]:/�`�_�MM�c�����Ơ���O��۲r0j��*��o��xԸ���Ek�8����������a���9�h����zf ��O���e�/�_��x�څ��\��M�����۵6�g,�o��D���Y�:��l��
��@>����5�'o�`�����s%Eo�6U ���'l#��P�?2(1;�>�:�ꇵ��P�/E"wIF
C��}�q��-�'XZ{����]�B2��.}�H��w8�^Q52��X�µ��d`�N	��	�.6+��G�&Ne���`�n�㮾�W⋛���C�#��C(����s�hPA���~{Ku^�lZv��t��ɪD2�L����;h�G���eCw��e_�*��􏆃Ӵ3���vJ�G�Hٺڝ���Gf�K�����8GWv:2�$�J�D��D�?�Ce
.�|���=�d�<x�9�;��xcߋ��t�����_�1]e1���c�K��G�1J�EJ6���������|�z�Y�U����܋�"���p�M�l&T��i?b����\z��Fι�e�u������� ֕Y*��(��8m?��Z�QcO����Gn�.W�$H�%�W��"��Z*�a|�(�9?G(1s�SM��6�,��b�t�����R0�nN�IX�%��<�Tr�V+L$��r�T�����?ـ���4s	V��&8OX�f~�U��/���\��D j1����Wi����Cځ�Xf�r��gҳ�b���u��{�V�f�'�}�PD�bF����(��;u�j�u�>�Mn�H4|�t�pme*R�v��q��276(t
2#uN�&5Ч�������ƹX�1�{��6�J�����*y��m*�0;X�H�XK�?ܬ�3����n`v��ᙗL�m�>9;��F��n$�]��qS�/�F[���qWr��,,��D��eq�a�r%O�$~2�@�w��SL3'K�k�|�z�7�\�R�[�	��	l?�2�QuY#�����,����`�:jb�;�v��h�
����z�\	V�i� �颱c%�	��0��}��9���n�Op�
�F*��G�f�4��F;
���g��ma�im���~[�!R�M�.Q�7��dd`�$8}ڡ�@LCO&�G��:�
���s%��޹z:��o���]7���� $G���2[�-5��?��M�����Q�g���2B�?b�����;zF�~�X�w?^�'�$�դ��ݠk�  ^X�;�����f�������*O��Y啭 ٖ�|���m��z�,SFp+|&������3��L�X+����$5�c���ԄT�_�e�%OZ�8|*f*�R�	+|���:)C_�I�u���$�����$��TN#����p��|�����3NN����C$��`����� ���;>or=�9l�vj��Xα�W��������yS:Y����F>p/2�t��) m�9�M�E�͋>oR|e$U��ϖy@��O�Uf����"8#�Bj��WM)�JE�t��#�z���^��F�2��
��јR��=1�
�"�}�@1�n�=�+m�w����Z-M0��kCJx���M��\iF�5�ꇙ�/����;��)R��M�*��9�0:Q�� �{H
(iz#:h����7`�p#'J��t�WY2&��7_=�W4�D��j��3/��:�#K�ߔU��y0P8kT��B��u��X7��~X���Uʌ; ��g����l��%H�(��!�����{�x�7;b���{�Em��?���FP���d�����"w sK�$E�k+2d�����r���eR-�1.��W8�$�7������1W
?���O�};���l�Lە7H��ƽ�0R|�T�:,Ib��MXj���]
�-�pWdS�P��0t#h����lo��d�S�` '��7���%�w}�cE�����Af�P����߇d����Z����lk�ˍ�,�}����oN�kH|M���#j��Q�Wj���I��6�9���7�7=P3�[ߴ�4����lK���p�wd��h�FO�T�J���(ю"J:������o��q��Ą��3)��r�=���7n a�ˁwG��&���XD_�U�@'JЋ��q�"o�1K�:G�"QlC�ә�X1gԀ�2����9+\o��8~��p|t�]ʺ���;��;�n�j����X@?�k���
)f�2r)�4��)Rz<��q����&w����n��(�RcNO�)�
�J̢ǿ���҄��f`F:Zb2��;6�� =UF��B1�Z	��by<\�_|�v�����e<*�aF�*1� [hg�A��[]=�[wT��yFH��KD.~�����ː�T6�z��N�/x�T&HL�p��T���B_�_�H�,m��c ������)�,2� W�F�$(�Msqv�`�FX+��g��r��W#��-��l���eK|m�&5�PF)Ք�'��8ad��6����TZ�+*��>�ci�G�:v���M_\�xX��xɗg.�ZH������Q!�c8`3��C�X⏬p���&l��>U��tyDX��],�r�i�1ܓ�Ir�*T;��)�,8����>���f����Ƚ���X%o��a��2D�T(�Xj�X[>,��*�[br���3�l�q�!����p��&z���܊	��a�O7^O�[sJ�.c�b�v0�l�[��՜�M؊�ˆ�`��^�����*����j�{��H�,��D kh>ҢD�[�RM�6['��wt���9k��������8�r�ֳ�(J��V	�Qo�U�r���]V���Z\�
:�0�v�/�);-A�@���ԅ8C��.��Ę������ӽ0��b�`�<%DSrXÒ'�/�@V5�q,ΉҬ����:��7�P�����ڸzTcs�0C�#tuc{X\�fZU���y��q5"VI�레_�����dSBryq�L�K����It�Wj'��P : ;�Dӝ10���9�q]�\k@}��	Q�84����X)N�.Gl#/�=�\��?@�6�gp��d^1���A�C��	��d��I���̴�
Q
VQ�-~s���*�s�
!�T,���E�4b�����{��I.I�i��� A���ђ,�Sx(�z�[G�����`� Wj�KB���&��(+�h� ���#�t(��f���Na��{��7� ��E_8+��� �ٰ��Ax�^�/�20�P���"5��!�����<t���B:���!��mY�9m�.�k��X0��YÁn&R�ꗶ.���2�B>��N�����$4-�ꔇH��d���W�����l���K�&�/�x4N����u(�Ɛ��`ZT����Nb���`����>�ZD5��8|�}͚��6`��>�=dȁt���=ѵH/�q�s��e*�fS��V���\�A����p�AU�e���,��'��O�w�֍~^cq��2:'G���뮴��[?�q���G��H���p���B���HurS���t�n�� �b��9��ή}���^�T�/3�qT�o6���&����k�A��컡�T+�VA���^��դ-]� B�2�WNN���.Ӿ��iE]w��J�u\/��ͅ�`��@�ܷ!7\���a#���O� �t������&��L����ڻV�L�� �"w�Ǐ�V��o����������^m���L:q�� 5X�/®R���W�K��M0�pJ�k^��:Cr'�^���b��dĝކE��ל�X��NP5���#�{n6���{ ҉�U��W�o��m��#���AƁn��7������w@�.�V��9�._���.lm�{�[𒪷˖�X;�5r'�c�Hx7�塛*=q=&~8�8*aH�v�l�k�}=w�@��G�1Nɢ|����9��L
I����oҽ��Ch*���^�������[�&Qq�j͵!�G��# �t?��U�ɋ�Z�V�� ��i'ǵ����*���}`
�_8y�� �m^�R��ؚ*%7�a��g����z��T*���0��wx�h�=��?7ŤO�=��$X`�څa���|B�O��@�xx��5����$
�h�`�M����$y�ҬP8!e�y1P�����s�Wէ�Ď��o-E63S?�X��Hx��H�����5)�_��J �~�G��S��������rU�L���A\�Tĝ��1b$�� )��ȍ0�j:jK�]RH)W�U��37�p����t�\��[�(���7�l�B.�x���@(+�KG�m�$N+0�'�wZ�ġC[�����`\ �j$�
�%f#�M��;T��
V0mG����@=�9���g���'t�����'vp	�.�o�KY8�[3�U�g��m�� =<�8������x�q��o9���8W��+ile��5��l8o�(PSi̾�U��I�y���>���?��gfH�`]��`�+�i�w2O�jI�Ѥ(v�¹�C]g���k��.����6�y!�M�o�3����()��*>	'�h�z��^��xS��-�8���K�Eg����>�Y?p��G���`�5�"�����W��ʼ��.py��PƵ��)6e�)ܿ�sG.֔q> !�6���}7��n������-,�����|�.jCV�RC� ��ǫ�HLC5j��o�-�Hp���R�@Ldc,��qt��P���/$']�P�N(N�A��H2�T����X(�:R3:���O���}�����dٍU8�J^Z���
�L�	��l�����*??����7q!`����Xh��|����=���W���&g�9�e�8���*E=x�&
�z������l��)��'���@	:��g��lwUw��G�53�e��nʱL+�n�C�_��iO��w7�o���W���=�g[�Z������*����@�t�z]��0C�:�+�g��H�V�PQ}�����?��\����J=��gh����/���M�Ia^��Y��q�@U~����r^�As��~jN�P�����|tu��7+�� �w[�*�-�����xx�͈�3z��ɴ�5�����kU��ŏR^�F�L{�c
4U��c���OAi���V�!!H���G�/s
ط,�ɖ<��2��b���|�y��ӼD�S�T�@f��1�aЊ�ު�b�U-���WI��ԽQ+?��#�/���nn�J������O\?ޒ��]bAP[�'c,��;L�/k5��j��#\�Y瀭�} iY�o� ���"�L�u�F�C�$�$IO�+��/x���`xSK<�
��᮲_mp��q�5�"����{Q7(���>5����seRc��1��9�Y���rg��A���_�,$t���`�[G�|�4���p�Ci~�nv��|:N{��L�`��H�x�����k���ϕ�+�֖�ퟁN����r;5�p��H(�#�6�t6�Z������mRH��8~F��/��?�CQ$t���࿢ٞ	=�ѕ b���+��Hb�p�#Ǌc
��c��Z���3U�o���J��q��8�����1@��w�P;�6��#"q�3j[�l^�%�A�`���Z�I����09��>hL�L^��G�^�clԵ�d��Մ�_v��H��y��� P�n�"���(f�Y��O/1�$�G������� �M���9���x�n���Z��޽�,�v�+����P������ӀS��H�H[W��[C@|����-���C�Ct
�am�QP�2t��=m��(���+-\�/-��@����g�t�m_I�X�YR1�F�L�ԂU��� ��㞆� )�8���l\G9�u|G� R��AOR�r/[W��k�k[��Ӌo�%��k�J
������Ԍ�isE�ɆQC!�� #6c�.0��<(�)&2N�i\�����Cq3�槦�I�S�ح���P��u��1�Jv^F�4!���,O
MffL$�6����y���j=;Ö.кN��
����2C��u�%�9�F�����2٠v��b���\�b&]2]���/*B��uu���j����k����S�~ %Iw�Mɺ?��|�V�{~Htr]2�7�dJ?�%��H� 1}�w`�����D�f΍a>����@O�O���"'l&B|v��b�0�8�9-{����.��پ�ϰZ�(��:
'����n<6��-[:�҆xP�I���q�-�Ђ<�4�]H�a-��Y \�y\�C|T<�V���m��g\Io_��3��)�K+�)U�H���sĒ�yD��k�zZ�����T�w�w���"�s���jo���kuF�Ic���֜i'F�%���1L��8LC'���j�����r<�������/����,/�;,�a�C��������Z�0���jG5�Kt�Z;�|�N�oL�ry8hM�8���i����-�!y��x$����(��;S���� ������-��BK5�k�(�9}���-��8�+	E�n��zj�;#������#���h���i]90�jxD�a��L��8���0� ��5*�q�*X�,�due:�D�'٣K���r8����f&YA[��'Wq7`4�]�D3���,B����5��i�?j�8���4z��W]�T�ә�#7yd��7�ũ\fgd<���%~�ܖ���=��.ҩ�W!Ğ0�G����Y7k�lY�elk8ײ��Öfە�R���nwTZA�����
�b� B+���1Ļqf���x�>�c���u��K�T��)Ggӫ2��c��|͒i��o�?�/	<�T{�L�Ј��y���>K�YQ��4H�csG^�H[������v�V*������%��Q3|.'w%Ƃ�4BiV���0p!�gL��+�����2	��<��i�E��,K��Cóq��GE֡on�z��w$_������Ի�(pǳJ4�-�����s�� ��r5���F��%����l�pe���@�1��UB2Q�d��Fɖ���ƓR�=W�a�(��#��]��p�>_VT�eIG}@�Y��<�j��r�%���>��Tb�ׂ ���Ӽ��}Ou5w���i�]�.��6��p"M�c݈%'�@�<!ߺK?��M=+�,����4���PѶ��N���?kހ��׿�$:A���pmW'�)Q����Z4���,�h�%䦞�*�A2`Z#��v�zOn�]�ɉ��tZa���������������չ9(k{"��oB=�a4 ���&
7{=���Q�����OBQ��fMDkX���#-�T�'���]��o�AF�@^���<���
��G!��7T����=h�v{BO�S����jA%�i�*}tVye����P˵���M5'�����\�V�?E�a�ee )��ꚤ�W��B�%1�N趺�:���wb��?�����3����[N���f̜0j.}`	�N�j��8۲T=�����:}���j�>����#
"�y�a-�Tɹ��B�R������3[�aS��-Gc�0[��Ё�oY'p��=�h\�՞�u���N�U^c���h[]����N	-\����鼽{�D�.&�@{@A�+,�^Bb=�Ľ�%�}��C�I�)�L�fՍ���F����_�r�k��xQo���	D��;5���ϧb6�G���ne��QCYer�m�Єh�wT?ď�E��M!�� �dE˼m	��U�8 �k^����X�/wb&���]��% ,�X�n�Łt�m���QX��C�t�s�G�M:~	6W�|"(,�~X^��O����l7eB����z��.,��ɔ��}Z�����_U���i�t���#SZ�	�¡H2l5��w�_�#�G�r&�^�� ��6�Ŋ��F3�L�0���,��ue_�r�{-���)��}9Rl
��($~(����SbQ=l��9�g��U�X�m�.��c[ ���7��fО=^�u�v�6C@���nJ,�8����00�����#!��d���]�5�F*e�T��훼Z���\2�S�Yc���Q=��rq�?͠�/�vE�8�(|�b�_��e�����"H9G��'F��3�yқ�u�=�Y�=�4~0������������ω�m�Im�����S2�Au����T5Y|m��l�&�xM��K���壡��A�|���)!�,g2����d�1#�|�� xH�N����� a���p��:�Ͱ~�D\��ޡI��Os��	�ɋ��ڂ �@Ky�6�_��Z�w#����9O=��q��*Xf�:tpeFb=�v��R&�����(h�Q�T&/��&!CPr��{����^�Ҥ�J���|M�\V�R�D����%��m_@�P�5Q���~��k*r�k��P����C?�f��$kq�5k�Վ�����0��k=I)�}�ԫA1#�Y�т�|�#}���i��'7)3������ki�-|��^�l�y&�ys��!���(��T��A3�PZ<}���}9T�$)J�ŋ�]8�Uhv7�g�:���q���%�LyK8�0P�QFy�\����*��J'��2���9 ��K�s_����3�T�zi�ȹ)�)�ov�l�ek�@�����1�#�Oj�/1��vߡ��="��oѝ��A�:nz21���X�w2E���z�ƀ��9��.���yld���%�Jb�!)D1Z���>Rr�Z��}.�j���S��ێ
���N���Fya�6�ݜ��q�il��Ct���!�	a	N�ﯗR}�O:x��ڣE��g�^��A���ge{y������֍n`�����0�6�I&�
tx4�	2=� )Q˫p��/^8*-��T6�C�D�a{9��:|N���*] ��Q�	��˖;��w��s��i��ғ�[Vau�2�K���sh<}�]؉�H���X{Hu~��\��g�8��A�:���Շ�]�k�346�gL[�B?	F�i�Z��z���a�#����qs]qbݼT%ׄ��*3�ե�}mx�4��x'�:�����Xy�g�>�������m^^jk��"�n/1�^���V4'l���6#��y�U$ɏ7���dv��x
��[����U�XQ�Ό7L|6�g%Y|�o��;�e�4�7�%�h%^���諍dm?r��߯��	�u2������5�������jE������Ezlj�%o�����|߄�_����bv���-���0%VY���\��p�V�H�#tN��jalg�O��G��Z�����f��@�#!��k���g`���#W���f�g��{b��7��1�*���y�^�p��I�7���7eMG���H(�(腳$r���eˣ`�v8_�5z=n��r�Q����b����u���~�#��Gh@su?���%���ָۛ�9\mU�2ȊZ\��ϭ����}Yl����w����,q��) ?����e�&bL�`����f��K�iyR%�)��b��ٽ��]�|�/�J�a��j�����]�*2�[dvx:4��h���1�ђ���kMs��FK�_�sg��-�i޽	}|X���� d�9+zü�裂qƽ�	]��E���Q�B�U����л�"ρ`׍P�#79ْ@����_N�S�L�>@C2��g��o]��1��>���3NYRK0�g�vަn��K�1c�X��i8�ϔ��]Ѧ_�D8p��?��iP�2�[͡EN�q��?�tM��n����X�WK��51����[�o��Eo��v^�P���Ժ-*n]L
	�@>g�[����q�N��CkG��M�I���f� ^�s�	�e���[(%���}e	5Yr�����B�k��~4�57�i�<!g�{1 �Eٳ�Ixz��֕6��ɲ.g�+c�xw�^7|�K�R'V2-�՘%C���}���sδ[�1�e4�ţ�x���!k�W�S� �������r�R\�I��=Qs��|*S�����V��u�1���A�TZ����|�m�J�D~��]��b�NaQ�I���;��<P�Ha1}�n���M�؟��|P G^��R@dV�#p ĉt��R�13b�r!����x��dŮg�Ƹ޶v��[[6�^�]E����F���Q�t�e)8��K��G�9�Uó���%�A	L��KB��ukx"*ħ�,����f�-��<��3b~�r�$DE}��lB��AA=������.#4-�ں�^���e�Iry�v���f"�aov�<<��ϸ������'���/t/|��,N�\!y@��v��8���*�����ǕXډ&s��m2��������\�4ҩ1�"L1u���W�O�Y�(Z�D�V?����*-���3wy�ӺyvhgPr��Ȑ��p�M��\zZ�L~�Qݺϳ�n�p|�Ӡ�&~d-���՚�G�g�<�B�yV�H�ш��[��I���3�V�I��^l�'��Jv'*�ء#_3������H�Q[����vE~.�l��	���}��Q��y
4d�OA 4ݝ�����(,_��A���|�%(���ݿņ�jv&)�g����!�����q�rT��ʷ�oM�>Z�(Ky���a-۲�>&�1HR�P��r�����!?��1(Ѥ�ؖc#ax:�J�Պ���yh�a���9}M���g�l�"%�޴��Q@ň�3��9F.������8��7�A�~�|�,��yV�S߳vH\�V�[����%F'��˹��[\��}H��^1J)��*�C{�9*�~ͽ�8���"8�C ̧=�%�TH8t�@�ڪ������$�V��5" 5�)zi��^���e�nu|��)}e� �f��!%�Q	��@��ҥ {+���j�*P^�h����{Z�)~~^nͲI��f����x�XV�7
�����N�n38fnUՕ]֬Q�q�TC,�w�M��X2�@�\A\r����^����2�I��
�70y�=�e���;Ss��C��\�������)�5V
sǨA��{�+�h=�*�K�2���#�Q;T�CZ!�t�S��J��}�k	e�P��iv2'XG���xcqss��K ]���e/���
	tڪ!��V�q��,��B ��q�6Qq�u��
��A�<���%�=�V(�}WZb!1��8քKG��6'S~E��:d�@�C�^
 �d_.c�`�gH�0Zw�5�DM�*8�'v׆5�h���~C;;&2+<9T����5>���d�Ạ5�X]Oa��ͷ�t����0u�K~D�!d����K�~b0���8hF��%��	�d
d�v�>�yߵ��.UW.� ���P�}8�=G����0䊜 ߕ�m4"z��8�bЫ�:'���%'U�u�Jv'N�#�ea���
v">�ߍ
�L����2zֈ'�ش�B�ύA��D^m=V���|��@q�Ɖ�������i`d�d�X׀���E#hM��:AX�N~;�&�
���N�}�=��S�_R����D��b��fk�F�t���
:��wi����%ּ�:���U[+{�A�����bZ�H/U
�g�zL:u���4��_��a�C[���Yn߱��p��%�%&ha��N�����M�
+�U��*r�9 Q�?��Ih���&P���{%!k6����7��QP$�L%oW���~2�a�����ᢱ�~4^���A�9ǜ��_�~be6�y��.���+G6����q�Y��4�����q*_��.�LT�;���"�}M�4_��ɼq�?��H�;8Hg;$!�D,�v�S�{�Ӑg,Z��e�N��~�е��ā���Z�!��(�a��LE"THc&f�7��ܦvs���iR�?�U}�V5��2���§��6�S��r�H[�U.���C�C>������i&v�F; ��t��"���K����n�������r#��L��A4C<Lp�˃��̷
���?�i�V��H2�3,BA�/���}�?[��1�rV����52���ϟ|�v���<�"��tb�x>��'�]�H��ְ�a����|���3�p�\'�,0��#�6X�EŝZ�H6G\%�Uwhz��6�
?��d-�R��h�QS�0�&��l�����}��=P
BNI�a��[����S��*Jg�l��ИJm�O屸���B��UQ������U�P3� ώ�9
5��ִ]շ,ꯔ�5C3yL�������TC����K4iP��E���-
S]���(<]�J�\�M���ě`���5%p��HKn���U�8@K4�h��Vf��
~o�|��>zE��|jT�Ou������ċ\O�ˬ�"���Y��-����>�M�2�gI���)q�Y��%�< Wv���p��ֵ��rx�(;+:ɉ�$M%����P�r1���&lս$A��g)������P�i8���{�^����/��Fe��Kʺ�n<f�������X$<�ZYk�'�%|)cc��qʟ{#��,b@�mꟋqڜON�[9���@�
�y���,�9��\���c������a�kj���#�tRZ8�2@!�D]�<M�ݔJ*���M1"A�Zp��(!��g���1rG�t̵*~�~��U]��'�C%2� �ѶS.���N��W ������;�`�s����w�Y哽��Q�)U�[�&g��@�#�B���u-��ɉ�sY0�u���k�]���u\0/�E&�r��M��\���U�����eZP;Y��Z
v��\�
�N�V_9�S�;gJ-�����r�WS�yb��c�.�pZ&\�U������	H��`��4�JA��WB�����A=$�hV�z���m�9�_��
��L�����$��-�ؤc����0o���!x���l�K��z �!���q��~��ϳ�h>��W#?GG��2�y�3v��b{���Qo����6"��.
d�2�c��(p�صſs�8���,c?v�dƧ-�*�m�+.W�Ҕ�@�C��>M��g��_q��K�Q�Oab!$�O(�w?�}��|�����_lE>{z�Ln��j���
�XxT�����x*�0�1Ti���v
��' ZOG�ڝ�'6���.�Յ�C�O
c��.���u�ȇ�+5et�P��lp�Y�.m:7j3�߈�xO�Ow{�4�r7���,g%����	�E��[�8�̉�G�6� �w��I��2��~-"]��~\0T�,`@�Os����?ck�K==�Ra�,��p�T�L��'��iA���DtWCc�d�R
�h�D��4.)�l|z���Tt�HzS5�"�Аh���%R�ٻv�;)/f�u��Á��v9|��b����I��o��[����F��k����~C}����	<�(�xz&\�}��!�̪���h sP����Ơ��:��tOx���'yW-3����{�� I۴抜��v����	��6��j"�1q�%Ӹ�y�O��V�aF���yL�V�})͞KU�F��2ۇ��:���K}����#ɘ���7.����d6巴κy��w��G�IOr���>􅴻����7�����������7�2��3jˋ8a�6�e�f�.��tD���;�Wt�W݁I��y;�$��~m:��sO�h�[�zgDX���"�آ�fr*�|4h�A��b��9|�N_�#b���IÕ�X�9�[r���]$_�a��.�;�	��sQ�g�u�	*�lŞ�Ґ�6�g	�J�Y�p,�ٲ$���o�ic
�Gjv��(8>�%���tb=Xy�W�%#�x8�4i���{O.�U��v�ޱ@���� ������9�I�Sl��W��6��#�0����2�5V1��&:2rɊ�}����Y�g�
}sA}�����Ow�{���"�V}xmk]V@��p�u�&�ɷ��JW��_N�n�K����v���,�ї@�l��/�����W��@Ky͝k�4�4X�N���������5��Wg�R6{��$��7"P�D�`��x�&���I���z�!	[�/\>{ߩ�U/���*����G����R��+o�
� f{����u��sQ(V8�|u��v�����v8�P��:2�!茭v*K�7��*|w���O3ͯ|Y|�2|+��N��3��w�%�&��RH�b��&��Z-�TF��$�u]�C�[��oi�ʭa���i���b����<����m�*/g}������	r�wR�[R�� w��=���%��S`�<#-���e/s���jL�p�˫�%[B�[�n��2�$��� N7P����p����f^��Ǟ����ĩ0�1�D?>�z�
xE:���e(Jy��'G�Ә6�H&
?2������|Xp$�.���Ƀ�:��Y��ӋQ,���]�%�M�IeʖzF�	v�gүO@��;Y�_m-=p�����]u͵��x)��\6�wn��'��*/�f�h t�C�J_�{tSj���QN�w��d�y���<�����t�;>�}�uf�Twphkx#6���E<�C���6�v�����5�����<+^��f^02Mn¾0ʯ8ފ��_������M��KQ[_I)���|	e�d�/����'V%���s]M/J��f1��e��Zei(]j8	tUoNn�-rC&�8����%�l���Q�;��G���{M�5���/v��i�{��T�,K�et�Će��q���s,Y���H<h��41����p��t��ك���Ғ�t�(#�r5gE�t�Ϊk�n6�3цrJ�O�m���|��'�]��3��#��#���ɵ��KmH����~� ���-���|��J�z-��?�X��#Q.�A߉�>j0�Ow��$�y��[��:[�N�<���~�.1&��/�M&��<�P��7��//u���@�|�d.�vu����&c�:��TUG(�Ek�ͱ�Ry���F���%��d6�=O8^�zE�!�O���Cp(�-��/�Z��r^u�Q�p`�=}��l���q��0RrS(�\ٺƋy�E���3ڵ�].��~�=xų�yG'��"t�P�j�͒�@j�+�����Y�ݗ=��"��=�;$-	���y²W�Ad�e�\t�T絰l���4�_�f( ��MݨV�$+v���JA�-���df�'.����H��*��gް���Hp�&�)���?Y�bf~Y�Q	Z�m���T �M/=��O*��N�iv���{�Lu��%����e _v�.��n����b�^8������K7�a_P{��ԭ�e��Qt��7H�n���!n�z���I=�|�
�3��;Bm��=華�_EL7�m��∿���� �q���8[��������)������H_���Y���i)	�#��gW��<�'���b�#�S�M3t�@��w���7�����̗p�m��E����S���;�ܷK:�u�P$#�Z��|�K}��r�¿[�T�3�/`�X�r�$`�o��Gy~DjyY�+dζ�<R����������Z���S��V	s\ڦ���i��6��� �8z��#g�,��G�oaoS�8��^�^i�m���x�;�#�pg
%�}>C���u�1�+b�=�V�����
�z$�ee�����YJ���y������A߲���{'�M�X�:��]AQ�M�#�-!�P��l�y����j�����S
��xm�!��^���`�l(�Y�h����'���㘪T,�f~��\Y�B�9��'6}��8�������߇�`�t8l���9���	;���|����㍩��6�2��,c���R���1�G���������[S��(KVv)ow����-�*�3i��V�$�1�8�n�A�q�i�U�E �uI������]�2�E�YwS�6ҮH�0���j�����t�����q�:wғQ�(��ogxz�O�R!��Z3)\��ҵ�_n^#'8�F����<ν6�c�/ֈ�נN��;#-��`�:˱i��D���^��*�nS��.�l~�tL		ۡػ�ml�/��:���2�(+�)�:��y4z����[fQ����o)t\���N�F��`��
�>���l�d֩Dq
!��`e��W���	j,#]���P���y{�@�N�G��e,CJ.�u�=��VO�\���&�8���%�8�z$��sJG��� �ן��#�8P�,�ĵ�)^�+����6���c�@��y;��)z�D^�6���ޠ�K>�y�7 ����8\}HE�#Kq����3�/ѫ^+xK�u��,f���ڀ��;���tx�۴oZ�WԽV�1!-\�l��3bSO���rq�cW�굩�g])�?��j�����K����׭'ⷹL����Ic���+��V!D�꒝��T��=�^Г��=?����
7�)ľ?`|cA�ex�/=5Q�\��kt$uǃ�kմ��{N2��������g  QJ��1�� �->��ܔ�{��U��+ꕒ�������j(�(�:4��J����N��b �pt�[
�$U��D�t��m.A _��l����W�5���|�
�3�:��0r��q�����
���Q�̊_,6Y2Y��v���v��>A.���M5��_�Azylk*˼�`���i����qOau2�LD�R��{_����3�r l���~�-�� ����W�y��Q��.��ߩf���~R[ln0w�����N
�Y��85Y�T=*]%���P��v!1"
���|�3�6|-M����K�^�������__ʫ��~nr#|o΅s.s:Č[2�&բ��N(x����H��q�-7@*�<cjrB�z��e,�R|����\�f������.��J'ܩ�gG���*"��ek�����$al�#�6@¾{��@�J�8�w	U�?����T�w�8��
ơ��"S�]���޵Vڷ*��8��̄4׫��ŝ�ͻ�r�n`�"S��A������HZ��C�*;w�OC΢u���Z��qY���G]�#�kK��ZŖ%�,}���wWád2�ᰨ��T���}v/��;��6�D�[����#^�Ç��4��i���M��4�6b��A,(�¢1�5q@[�ߑ�H	�qs?CdH��3�E9��8�5�8�/|��aߪ[���r������I����
�/��ĭ>Ku�]ӷ�X��5�a��U�(K���%�z#E�x��Sپ�`�M\��^d���p�b`���,&Ăi�J��t!8WI��)�vM�τ�S�s	�G\_��-��ˠ!�6�	"���έ"��qB}���U
����ٹRo'�>�0Ŭ��4���G'C�>�U%xR�~��YEI:�����o�0�5
�h��4ǧ�B�ڮ}��;^i�d�0fx�s�u��H*B�ʒW$��\����������b{U�Z�%�'���w��/��r�7gys��c�������}~��ZA�k�"H��ӧ��=�|au�6Z�&Z��;�ko���L�*�+u���{LVU�F��q-4Ox��2����_���	�)�H�6�Md������Q��ڠ�����]��R�GN�
yK��UkWִ��f�;N�6t�� W�|r�7�C�.�*C�t$_ڨ�x1�⬈I�4e��ݬ?�kE�=�W��=}���'$DcJx^G�J�����T��7VG[�H�;Ǵ�3�|Y3�G)�S�a8�4����T��jNեenh"}��Aٴ�]�n�9smT?�r��2Y���m�4=0	���ԆI�"��Jp��"�P������]�M� x��`A���#�r�Vr�7X/����S����=V:J�la3�H9� ��AEei�ק���Pچ��OH�]�o'/�wN}%ۀA�X&Lf��9�K��2��6x\�
˽��CF���ag���ĂK9OׯfAִ�U��^l�����I8b���_������~���	/�r�A�#:�MA�~q�XE>�4���c�I�^T}�sZ��en�`B���x���=�El^���^��XFG\Y��`�<����2�#�Ēs�',n"t�R��x������ϟ��S;R�wG�Q)~���S?�<��T����v%��W���x/�/	F��p��.1r��=4�j.�;�ݬ��O
p�r0q�X~ FeVQ8/J�v�%�zRCd9�'����:� �h5Ƕ;��	$�;�(a���*�
u�%E`ߛ�u���8QT�:��R0.����Ѧ�E��r仝{�0�!�'W�����A�I
	�32|�"�G�A��ԻW��!
�f�ܝ�����+A�'�~!�����+}25���u�U�OU}VU|:v� +KQe�!;yQ��\o�%%��" �������7-~��̚�nsc$���������[^/��������|�8h���Bd��~����%"*��#9��� -_E�M����=Ǐ�k�-���pu�M=)�t�f��'L臕SO����-�D>(LD�HK�r&�z��S���j�~v0{��?C�.^w3��E�ʡ��K����,K�R?�G��.vc��ek}o���XeȆ��j�B�+��繭z���Q@+��O2��.Xlr5��2&� f�Y*Z�#�ٌ~���G�f��W-+���N�	&P4]�5q�<'v(l:�lS���+L��<X1�F���G8%I+?���}�@�V2�ڔ*�mR��	�]։!`��;�8���$3�b�J����[ :~B�R��K��B��y���<�ҏf !/��I��ڐg{i�����%ӭ���;��U��d�������>1[�K����r�'P*/`�f�������ƌ�k!B��=�,̿�W���d���?�����a�lt���?�c�|7�uT���).� �r>��)y�!��ֵ�rzM�vp�Hh�`���gH]R���s
SF��G�Jp?��	)'�� �;�b�'�>5�v��c*�'FH�@N&�m4�>�F�奕 t� ��~2`DMZ�Gu�W%���b75 KH,}���o���� ہ)�Dr�;\�n[)�jk2g��cH_�~8%I��ueu����8�*��t�����Ko)��[	����$8��1%�^��������U�	G�+�BwPs�׏K��FF����'�D��W�h#����{������U�a�Г�K倝:�4Ћ�Q�>�|�c$.�����/u8t�>��x�B�
J�����<��9=�[\蝯�)��X������Ç�ń`	و�=��2=��#uV�kSW�,{���2�k�w֑3����'�8Z���N�����`�l4ɾ�hG�9�7�EP�y�������J��ڜ�X�o�����}�+�;�dns�
�'�}�y�LW�����U��r�$B��:��8��tT$�c�Ih�1��[��w��a��XM)�5zQ�M16�i�z^팈WZ���ߧ�RVL@��x��8I�pyB�9=�]�EV!�!���jR!��ҿ� �f �t��X�ٝsTX܌Þ��w#��%��x�HLH�M��+%����ү��Qn1�J榐�<�������?��P�Ros}�v蛿�.I�㒄��1tS��� ԥ��J�D�1��ӵZ��ŷ�Ix�"�`|���� a�h�R�W�����ψ�9\�T0��l�$����hcxeX�����5�_�	�XD���IٹmFP{0�[�x�����y���qD� ~c�����d>j{�F��v;X���<M���@���
�#�Z�q1�2��.��JW3`�$�j�
���[)��2[|����DO�m��Q���!���m��%"N�wf�n�[W������6H�NR��:bg�RP`7_ů#_.)����i5G>�w�ХH�Z��7�����ەl���6�~}��}>mm�P�����.����{·Z�B1Jd|tPů~��D�$��
��C
�����*�,`q]��O�(������]�|��~mI�H���p�Ai:�&tP�GjϧN|J���6&��$aM�ɟݟ��N3[�e�L�m]Q�O�
��?�;�¦ul�K��H��)����a�O��.h
�Ӈ��D���f	��V��ͺ6v	��Z�pzXgV$�/��{���H�Eo����㲖i�~�b��<��v��L�T�a�!v�b��U��jvus��ޓ�<qy���I�4�}D��4�u�k���9����UKb�v�l
��<%�7��"&�<w1	�[�#yڂ%-���!�ӻ�7���߰UZ�`6F�#ND2���������G�eG�s{��!wCο*��ݦ?��"��x��d8���[��e����J}�?-��!�<�j�`Y����"� )�C�E9�T��kY�����Q��z=Ȏ\�_��WjC��#�Y&��[�0��Du��8��Ir^ֳ�I�JVz(v�����J����}��cʢ� L��(�E�&d쀹i�ړ\�6��r�Ѐ�7�ʱ0�\i&S
\(�z���s��
͒��F5�[Q���H�S�#?Q7����g^�3�c1��dy?��u��Qv���5&�`0����;�'�U꟧s5��C?bWa0�O#0����m�o�r�q[��2ӫ��]�,�TZ���V~Glq�h�KV:ҁ ���"Y����<��N�l�G�r}�)`�}K���Ӆ��x��4�4�����Q+�S�� <�����N3ײ��φ�j?�� x�)p�Bu��k_?��3��$�ڎ�<C2�F�,���ލ�6"[��=�0f�TQ��t�:�J��(Yy�9<�G�J�A��5/#���tI��]��k>�X��!�g���Z9���56��s̰��ڹ]�3g��tt91�FZ��Y�"�H5�<�G�����qx@���'蔙����C����r�P?�{�>������H�_Q�q�vLR������d�xp�����%6"8Fq��C?7�5�"$ʃھo4�<��0��cׅ?�^O��9F�s}�O�BM����>�d��W�B�K/�鞟�/�T�=��З��a-���H�4��N��܋�>�?�>x8����y�F`��D_d�љ%=���^}�f�#}v2O�	40s=��:��w���'Lʀ�����Ί��������_	��kh��Cc����%�?_�íXN�[� �����!���Bi��2A��+7�=�������(p�T5�8�
:P�ޯ?tk���d{�R��%�)�}`�)��q��j�t�ʹ��qnA�	���L��L���� o�����U&�7�o�`�e�oǻJ�H�����'$G��f�����B�����%����܈��������U��J/-���BA����K���O�F)�D:��m���^ʊ���ڲ�T�q��4�%,�\��~����q����^{P�D�@[�ˁ�@�T�" ���J�*+�)U`����`��97��rD����.)���tC�]�Y�ԃ@���D{�����&|
7���=�6Ǐb���bҞ���f ��We��4�:�W�h���z�f�5Jfem���AB�����:"��WD�u���_�����m�lB��g�Y�^�r�s���a��x.[UG��~�����#-�̏஠޲D�E �����3��/��zY��:�X��a�LIYj�p�y�3��iĞ�K�}�袢�S��O��aᙒNt�a�SW���+j�̐��E2X�8R�ں6��J��^&S[�H��u�U�u�o�f�
�x�g鰿�j9xRF�Qw��ŵ�ޓ��%"J�8+"}x��	-fD�|��������T���3�'sW	�~_��eGrR>������To�t��0I��!����V'h�߾�E���&�I
�g�Wyld. �	eN�W7AI�T����j���W���_0w�D:��=I�*����_�i
x{x���,��V]�v�Ӳc]��O��d���R��wlH��+=�@�nLyW����*mv?!m�wJe�n��BP�4��0�eݪ�A�;aF	ܪH�w?����䖯�TR���y܁�i($�u�R��h��l�4[��;���oA�*�3v.����z�F�H��B��Xg��#��\1��_ڳ�$��U=� �Z<Tȯ���z��OFZ~O�"�Fh?�8�p}��]�:!�!s��1�Y*UP{��{�w&�ۼJ�����;l'�߇� �y�����fO:H�޻~��|Y��u�ӈ�`h"�)]�{yG�&�	�/�E��"8)�䇢���{f!���tU�aؕ1�3G6�B��m���"���P�w�E�I-%�qI���F�:�A��!VJJ�Z��+,��� ����쾛���l�bK���c�P1J�?����yi,E(	ŕtr���zq�C�hl��m��E��˴2՟�СB�:����%4�1��2�����z��J�[��Ķ�t��`�[�n04��:)"T)Nv�55 yD޽D4lP�$Z&.�4��*`$Q�*Z�7�S�P\ȕZHM�3�u��������t�p�.�Ξ�_	e�F�L�7�͇�mR��u����A{� �j"�Ԡ�6
������\��%������2ϻ/�_�"�䱝Y@��������������Σ'�C�q
��v�)"@�E����6�D��;H6���k&!7�б����u=l��r��{�J�2[�4_������9���r�D`�;Ӆ���M���	���Pfu$�x���|h��|�^��}p�y1:A��"�W*��Vǘu�����cQj���zF��e��&�@�sp�Xh"�V&�t����D���L$}���d��tb!F�}��� �]O������@j���I�_o5{��\�V�N8;�]�k��Uh�I�!z��Õ�����t�v Dg����u$���|�����g|�p)�#y��"�ba��=��,�����H���-u�����a���Ǵc�����Fg�W�E@��9㭩�����x�Tpw$������<o�;��H��J4�
:�H[�҄�+�a�z��k�1��آ6VQ��̈�0���r�q�D��7<+'�;�X�V���:�W��tm<��6.�8u��f��J��j�8�zA�Q�nX���-��m�ƣ������_ �6~�9��� F�r��,܀�T�gy�5�������&�V~u 6�
O3���>�|�,8%�E�d��~m��naO�����.������(&,e���}��_�����>��G<3N~�E�aF��g��y�C�}3�����+��_�v!;������r�I��q�,��U�c�w�Вk4��=��:�ezL4 �P��?��I�B�g89� ٽŴY4 ��-��d´�~b�����>��w�9�u�	���׷vg� �F�~-�>�P��=�@c�8�X覜��fܙ��C
��
]H\զ�$���]k��.1�dw��Q�pB�`K�]���YEd�ޥ�����StМ0�@"�]���#���w(`G���*�T�2.�-O�{eM�"'ї�1�j�<\V�?VU�*K�*�[E��b�ը�O�U*�?v�W���fu�`f����� ���b}���(�O�t�UeA	ܝ4�	" J�h���%���Ti��k)O��|��;�����Xpzq�P��:�\O*�]X+A��]����br���)ͥ�2��~��iI����0hs�q�l>`�.j4RB&;��&Ia��#����^�|_���s����U����vVd?��\�cȬ�[�� #�i���N+��D����%0\�N��DP�i `��~��v�9c
��=�K��m��@E�w�pՏnk97d����E�z��?n�XŠ�m9�qUb�{��EMj�
.	��)��e���XTߐپPq��@-I���y-�
A2�������Y2�
�^!p�u5�ԗJ��1��D�	���ܝWw�#;zd��ơil� �>��f�ᡃ@����뽗kPT�ju���O�6�l�e_�8B�
7z��PN�� 
g�a������_��W��$�i�qab�Hj���z�I�#�^	�� 	�S���s�v�������b8	�m�*��y2�
fxt�W�vy�ג�� -pV5���X O5�ԧL������ԩ箒�n���g�ެ��W�\��S��-����DԀ�O��D�A�u屙��|�ʥ	U��!��?�ͅLY� ���H
"��H[��O�kI���x>���&k�n�p�_�C���{����h���wp5��ux�qV.K��:ƞ1V;�g�ؔ+P�!�>Sn�Hߑ1c@~�����w�<�L:�ň��Ag�F�d��71q����o�Ƶ'���E����bx�x�g�\)HUy�����ī0U);�J(����������!�+?DV7�Ŷg�+�V��� ���N����O�ⴚ'+��*�2� ݆���{E���1���o�O �8�^!��M�JǾP��a?��7��[�{�i���u]�b<d����l{P�c����'����u����O�Vfo� ��/y�������Diro�3*������lq��|���P��EQ�[��5.��˜�b1���ܯ�NE�M%*F�26?@�������|��zW��@fy;��5�����U��K���)Ŧf��/"���8E����B5E{�����/p�M5e��M�AL��N>{>�D1�6P�iPJ7���L4xG�߸����F ���M��z4�P����w��ӈu}κ��a�̶����;=;�'�1	���[oʻj^5*P�ѷ:5��O"�����a��y/�Bӎ�ш�ևF�xSa�y��^��&ݢ�#��1�����}Efǥzi���%)3$\(�$��BV4e���KS�`{�p���B��t��0�5�̹���V?2������$�޶���r9H:�q���ZZT誒m�K�޲�T�V�eJ�Y�0Xeґ��_`a2�U�{�t�?�� ����p��2�%�7�j�޳k.�ͥ5y�g;
��F8��ˬ=Y�,��
��Q�����$b (�BZ���0R�����ϲ��wCg�mΩ ���������|�R�x�������t�17���5e�K�-\�ObPh̏^o[O`�����鋿ܥE*_�s؈�	��������'�BC����Rs]�1��m`\���k����N��D��T3A?����!��-� Lk���Tu5�ݤd�-���OՀ7���%�\�3t�;���Ꮕ���@���I��IZ�v��I��B�H���8���N�ֶf���i����j�&�OD.yG���*_2*�zϓ-�+hFLi䢣���>�d���p;?��]�K��$�w�V�F&(�ݍpbwȅ�bw36��Ԏ���fZ��ƴs4�:)��c�@N�'�����"|���Z @����B0�/��H��?�O�Ć����D�gG_�u+ !ۤXɓY�>����i�Ǡ+�e�ùd� B(H�9��qHA�,M#/�T����&�]#Rd��Mh)�yJ���-n���(6Q�uĞ7����XNj���^��3_r$z
(�X+��v��O]�����dD��Sƚkt�w�j/nz�<Lk�(Ȝ���˩���l��qkޠ	3�J����zABV��y�ߍ�]��-�Α%�qJ���*YC%�x���}��}���\��N#yn�R@��_U:���@l�����z)��8��q�nkF�� �ܮvs;\rΰ1�0[��d��A�g�+���%����/�v��-�p0-����J�����;�駮�lLi�G��N��	��"��h�����8C�����t�
2Fr�����/�զΖ��]3��:˸z�r�b�)-Ί�����򮌠z �@yK|��r�kڍ`w����l6zDV�ʑs9�:X��T@Б��.��w��z��Pb�������[3�{T�wXR>�"���Ql��!�*� �$�S�,�������)v��)Aχ�ad� �M~��&�Q��<��f^�q���
U��\j-�B�ѧ^>e8�v��qj�yZE����oMl�P�7����׎0�N�1#?+�.�:k\ݒ,OЎ�<y_��р�V���xχ��Q��l�Z���Ɇ�ߏq��N�����G�X�y�2l�д����~�����tG��`���~��ذz�5_�ņ`�k[%��������E�L>Q�pFt�J�~4��'f/s\���-��L�r@(r�ķ���
.�(���Y�!���΅Ew�O��iu��rL�a��D�;Y{��*pn����=鱘�n�����wREV�Li���ǫ�FU4��� �;K^~���Eg��3��i�S���Ї�s�A~�7�.4,��s�Y�?;��`�1����v��D�s��>���,U�M^�7Sz� J.K=��pv��6j�"���o��J���w�4N }1�����g������U�>%���n:�_s����?�] u����\\����:o'�քW�����0��~ĕ����5f����(�
���g��IY ��I����ԍ��Ӧհ�)�H1�,�B�י�cqɤ�Əm���-^��Ex�/]��aј��g��CF������U�T!b�k
v���%��7�%8�e%?��i�I�d�@,][����Ü���1'�&�GG�$����ܽ����T���6���}����iШ�5o�
���Be�t��q�ߍ�!B$B��z�5��2��O^��X�:U���F�|OK�}�x���4i��íi)�V8�)��O��r���F2���(�y��I�93�:H��~�j�b"��f���İч�8���ױP[�����s�&�%�/XU�>�������ei�9:}����0��+��z�=�Z�F��MCw"\ct�8.i�2���}@C��Ծ��8<��j�����y)*�b�Pɱ�c�@�፳���<
�V20d<��c�����@��@,}s�B�''�	���)su���t&lP�@�����c����(ynڻƬ���7M�!����/�zj����`Ш\uV���tZ)e)��-|��˙'9rtEi�L�g��Mm�,��w�q"�?-��U���? �����V#����<.u.�d�B����xL�;h#��h�ދ�����8�#��|}���S��{��QXY���
�N�Yr�\���Bܕr��׹t�#�����h��P�k�I�|�|7�Q��%�Y%��?�������0��V(s�8�I��sxGz��A��Q�<4d��_�'|�Z߅c<�)-�/�+ 1$WE��,S��VA�o��P��6f�?(߹�R����2�8b���!?H�݃|������@�}s4�3��<w�UI.���>�HV�Խx��܊��#�z��I�����A��l�tF{#1�eb°���(�g�:�j��^�by�XX�h+��ʐ.���.��
W1�pu�KD�����G@���/,"%/"�B���t����|����t�:�˺z]t�|��ID�!����ɐ���<v�������c�)�)��!���K5��rʛ��$�/݄�8����r���Ӓ�z�Y;���@T�!<E׹pȷo��v��zۂ!�բ���K����r��90v��~�K�(��b�{��8#�E�F_��^���PQɋci��7�.�f����.5��U�m����.�	W���ix�l��<v+&�/W�7�ڑ�K ��q��Hb��=M��m��\���JjA��� f��Cz�з�N>�;�M��#✑�^�k�O;:��̈́�.j>OԆ�R�x�չ�8t� n�x�O!*�(tɘ.��)QC�q�%��ft9ܪ@IHɮ���{5��Ka1��틳v��Iy�\"�,�fj�azw�� YwTFu�?K~f�?�bS�M�]�\��Y��h~A�/J���Ϧ�ǆ!w2�mb�OܪK����c�5��n}<fjv~�q$��Z='��F�!����2t�j��]�rzp�Lr��qMʊ���ӷdM��?vD�H脏���q��/Ւ{��E��W]������Q�"G�A$����Md�}p�}hb��_��Հu�=�u^�m��r9D�}�+f��,w�����,���2��U䖨Έ�D�˟�*��;V�GV'cr"�`Yv���NѦa������џu$��~��N9� �4����_�V�+x�b������*�Y�����\�u�V>LV���Ft�a��? ��8}$z���sQY�̃�������?�{%�,�*/��1g��h�N�#׶��4���V�秡x!��G�\ר<���l- �b�ڼ�����J�X%9��?S��2�r&0'Uב�f�-ǆn_�LJ\0:qT����,���������KJ��G[-$��&dj-�d8I��5��=�zVL��X6%E+	��0�b� �W>�-UgשQ46��G���⌲�|�a��LX!r�Y�z�����l��n��O�����H�#����j��ڱY�])��"J�R�{�pW����^(�i4r�l�����;����<Gä�)�J4��k�\��v�j��X�0dR74�����3�4T��O�C>�ȉ�߽Ć#�\��M|��ͣ2�~�;��b�;0��1N�]�����=i��ӗd� ����%V��
x����W��2v�5��=8��/��x
�IᲣkB��7/����R�d�bW�r��c̬`㸄jIS�����z�B{�5�����?Sp����aN��t�C����z�J �o*�QX�1$@*;U,�t3��P��A����P�`�:Z���$�ӎ ���6�ˎhAHu�x�R��W�F��썭�g��B�;���'��ne��أ�B^w�`�>�E����d0� �u�;7E�kW@$�F5��ޡ�}�ω�S�|!л��M��L�������m�Ttۻn�"�}�^D��h"�����CH�V�nu��+5L���5p	����톫�?������4~Y�2v圙��2�k~�=6P��{�G��I�`c�'z�g�����nn��]�ɥ������&�I��p_�<>_�׶����J{㘧�B�2����J�1����żF����;�"I�_7��?)�/�a��p�u_>9���l��ʇ��r:	_r+�
)9N�.O�e_s��x �	��D%h��ɾ��o��@hB�M d�0[r\�7��젅�S��p��ز���Ժ2Ę5�Pܝ 	�h�V��b�9:OXs�1�_�N]�c+��-��I��ق[�{͚�=��uC�u/��F�]��l��Z��HH?���#d$"�A�6�����w�E.����TM�ƾ���]V�[�ܮ��D�{z�E�@9���u�~/-��HH�(�O{�����$�ZOJQ��Q^�q�[���p�EK&���f7�rيp䎣R���Ο-?�[H�{+J�K�c�ag��H��-����
�����Ƈy�Ew�_T�=;*B-jL���L������:Z[����\���4�0w���~2l�h!|O�1d�8XoR ���K��s�9ӭϩ͜N�W��5��Z��w�٤�n�nP��X����X��	�y��SU�J
� �Oa@$��x	��,{�4�F�s���½9,����"V��B8���Ӗ=][TL�3V�*��J�=�`��?������I�������Xޡ�v.D��r�a�di���y-y���K" Syl�� ��[�,M��И�7��<�2�� �i�d	U�d�������Fbw�o��8?���}���4���Wdms@aL�c��@2���{6�W�8ݕ�EiƃKGGxT��`�Y~�;^E"����tƏTK�ie���s@����/G��A�#��f&H��_)����GZ�d�Ԧ#���[�[ZcnU]B�Sf�x�W�v�3h��K��ڋ�F=�WI�Y��w���
��G���<�PZV�`���sD�\6�b��9�:ES�Y-c��bԏ�S���ˮ��"���*��V�a�olE�"	�!�9	�oj$\�@3�$� �pz��H�Ǳ '=��<���x7m|�B����T�?���)o��֮��9� �M*aN�;�>�:�����8re�ﰀ�ԩU�N�{�Ͼ�4jG�K?
�_6P��sY��n��ᡍ���E�1s���d�^���3�ˊ�f�'����D�t��ޅ�`�:��]ܺ����OWFl��.w����S�(ǭC�A�Ž�(�!�bd3��D����YjDo[�W������%�8���j��U3�W
e_�W��s`���R@VPY���jS9\�"��m�ґ�ic���4���k=��3Z˦���8Z.�3��u��LV2� e,�X��P�=D��:��R)�rP����-����L�����_�妸�.-7	l���3�W�b��g�,�+s���D��@�S����\�!�j|��R��X��ȴ������T+F�خK�x4KA�}�/�~R�M�C����~���s]��	�,�-R@�JGSw��-ywJʱ�au���/s�+��pz�?)�eqNL�ޢ� ��gx�2������-r-k��fP����jY��Lc�S��ڠMPu�Pit����1O�p���;�@�f��Aj�Z����������in���j�ϗ�| X��������]���ۅw�%�J�����e�˪/���X<B���}�*~6��z��& ?��T}%r	q��yɋ��)0�8�h��^U�NT�0�^������İ%��=rNw�ɦ3S�VU�m�RL�ju�T�y�k�_�mG���->�`�亂���قG�urŌ��/e�Ez�}��������V&���G����kȺA��)�!�[�ƿ3��sM�u���5B�6�dC0�)��CP�d��d���'�`;`��߁`�W�v*�c�f�^@��,�4f-S��؛���k�+��u�?�e �bH�r��^J������2:-?��Ό@�h�Q$��yr˄s5�SV缅k�cέ�hE[Ac�[r+]D���P��쩬�~f&��see]�)(�=C#� �}W�F������QOBN(d�S'������㔿s��ְ?�.?����6'���.�Q��z��������XZ�{.�e�u�ڽ#����BF�-�U��3�d(�K���������(M�.X_p@���U_!#������GC����*�0ZTgG*@�Pfo�U%$ Ѫ�B�}���&9U��s�H�u|��C��e(-�oq����4�j=	F��@G��Ҏ��W5k���Ȥ+ ��Ƹi4�@<�M���[M�r�.6�؝��9��O_��Zʆ�]�s�=߫�76|tEb��~��
ϝ�L�|rr�����t�6�4��?[�2x�k�ܔ�𜩁�"�1����ݕ�y4�ؽSE%3�d���ʵ���撀��%JM+!��X<0��9�ɷ����&�.ߩ~�����:L�m�[�z�ėU�e�d�1|�8f����Nn�뭳4�9G�:�PϘ,��뙀V���[8���M ���K[4���AHZ(��$u�CqfK
.������Ǐ+�H���6k����{揼xı�u=�P)�l��M���"-�i���a�
�a����77��#��b�,���Ft�d���	Y=Q���^�������*��Z��|7�%����dH�&���"���Lo��!.����ɂK䂒Y�"[�ȀڤE�lk-x�-�ZG@8�p�+�E�: ����3����˓�2F��o�!�^D$^�t:�[W���ԉ��÷�i��ŧ�l�'(Q�q���q\@�n�Ɲ�2��7�Qy�}_VtC�ы�x���"CM[
>/>|�2wU�ޫ1��ڋү��Jw�%��-nAK�(6��3����cN=Ոʌ��
� { h�k%?���W�}�U��3��b����]R�v8c�Je'M4���lJG]x���� ��f&�\L ?xL�Y|��nfE}�1֟��G7^���&W�aZ�C�m���	5%|9��?/X�R�V���@����<��?iO9�O��S�����8��q�Е�IQmƿD�=�qQXH�Ӻ=	W��6,�7�5������e� \d�E�(|E3�8=߆��H�%�n,�����{/��zϔ�|̚�=�o1V�_b�˼{��E���M��~�Nt!�O���ْ��OʍP)?�ɳ0�G��+�/N�Ƅa���	�Y��ۧ���?��ÇM�J��]�������:�J�Ŧ���&�ʳ ��`	�.��.nhwH��5�ƚ�@Xm:���#�͸�a����f�r�j�>���h��U !
�6�i��82ܖaۘ�u����GwW�2�������>͕[��"jn���!�3;
<�.���S���R��-M�hwh���N�?a���.�n�e��>�B[�`D�>@転ϱ�"c�b?����Ѵ�s5�}F�{@���������c��$��2�DzCJ]�4��H{x��ɋ i� ����fڗ "6�y����2q�U�Q��zl��0�ҕ��*�Ӗ��!���t�������ٝ�ǆ�νM�ja��l�3���Ǳ�?���.s9���G>p�E���Ɇ�rd"L�b���uI	����Π|��s:�R�Of� g�Ds�3?�U`u=g���Ѥ����.G0.�NT�P��峺�L�0��e��F�:�)���ՀL��<*#����"�o@��)��۟S���͟kv��,�!^"L�O	:3�����V���b��ؚ�3�^L�5�I��'D
Ո��d9-a{���m�K�M�y�j �iNJ|�(@$+�x����ߛ#����=jy"}�4�n\$x�B <8er�Α�F�:���9����E��nϿ�J�ȳD�-·DT.�yé/�K�Ik�l������le��s����$.�E�H�9,4w��7���G�=J^X�ʕ�_T��S���.q�UO���
�V�>��3��k�K���9`�<)�)���¢
KJ0-���}��a��� 6��mH���Qm{��(K�f��}^�E���]8�,BW;w���pN���@�:l��c�|={6�$$:�F�L���9TǪ%��8�6˿��@0��w��6��{5��9�A�'�R��q]:��Q�/�C��1�v˾�qg��[�[.ԕ@����v篦h��m��g���I8��k2}wH�W�,�{g��k����2X|��������z�஗���[43R�r��
�g�.��bf5cs��yݨ!d�R:������l�I!���2��U����$ �u�oP�8�2��7���׺����N��T_wz���(�[�����I�#�0��?*���/:n���x�!�p:􂡑j�2�s��K=���B�zz8�N���K��d4n�\����k7SBP�x#�i�8�j���FԔ� >�I�=՗�7�"٢�	l�n��4�bUy��g�a��z am��/,�ʝyN�
Z�\\���S�]x8�#&<���{!K7]�(yk��L�8�(�L��Ys��T�� F��])6t��o�W�gq-@X\U5c��b�@e:Złޡ
����̞{�M�; ��T��D��1�rq-�,���#�F��gO�<�0��6n�T�K��\���/������r�\>���8�ys�e�&?�-����;E���j����	|)�bg"�wң3�+�'}���Y��l�J�U�wfc�!>�ی�r�'N9�� �vRkO��ӗ���yp�y�L,���;<���lNǔF��$#6��p����n������w}x��$ϼ���&#�C�7�4 ����[`�b����ݶ�������������4I����.�&x��f����p�T��ˠ�b���s�m�������O��!P\�f��}(�ZŨ��gF���kQ���N:��C_V���6���0	>^w�
wf��fG�U��Z�l� �-��L�yų�PM��+h��A���ԇH��J�I%}sE�Px6���o�l$��R����,���;�����a�ty�4s�
ZL�{�����aסԬG#l(%�g�x"��f�L��he�s�`�b�!��������bZG��5����)�t�c�G6���>���d�K��`�faj�ˡdq^���Z�] �����k����Ј�I�P���3���{�>�S��ɋ[I\�:Ż2{�F��%~��X4*-	��g���tFY�<�(8��[��E33���� ����K���7�B�7G�[W;��|Ꮘ.�V�I��7fM�����i� ��3)��SHK:����O/9?<s�(ـ+[v�����B*U�^�����!�a(X����q/O�F��{�;C���V����l�5[AW��jh2�Js��ho*X-�^���C�W��T��1 �n��"���*�Ɠ�oz�FEK����fz��� ��g�P��s�DD��A�b�[ܱru}���  t�O(t1h���~�O�%�@�	��یo�.�����LSo(��{�����ڭ�s�q4�<���We7=�z��	tI���@�P�r_,y��٨N����c�O�߂0Tl쯜��`H�!�
�#��rRG0�Z!���z�g2]��|ʫ��� �e]�~y ��+�{�iu�8�C%m7!P���QX��=MR�_�f{ʩ�i�:i���6(�	s79�� �tJ)���N	C-#����-�>�漙wVY�G/CP�˖�D���S���>}��F
W㸶Q�9_�Ϥ����F�]�V%z)�\��UFAE����Z�¼�,F�9-�q�*8��C�"Z���B�A���d^��t�_s�K��/�d��V���e��柎YA������vz�)�x�s���}��IG�����MJ>Ko�ct���rs��alB�;(T��D�=�^���8�%�6J��:ĉ4�}=L^��ǋ+_����^��ŉe�j�>��A�篗y�ۅ	V79sI�LW�zu��Ҟ�3���H��C��t�e��Y��� ��t	\�L�Q�	��۷�a��� (D���T#K�K~7�%'��/#&m�ص9[���%Q3#������5�n�?�=7�4���%����{ɴ�2y�8��:��8O��&M�q��ݽ��;��c���[�M���.T��fI���+ט�V$l��ۜv��Un
���}�n���qO���"(i-q�5�,;�# f�"N��쓪���7�j���7������9��@���r!�<�^kX�!�09]�j�� �`'�w{�&k��\��"(B���N� �a��"�&~�̧��YfZ��e�?� U�	��:T�*%K�&�n�ݚ��� Z��B�s�Ȃ�;Ԭ��X���<�0�[�Ӷ�����'��8���l��"D�m����W��W)X(��f_��rw���]�&0N��8�~Sxf�Nr�SO�L�g�büp\$L���y�a���C������'�R|��t�[�J���_�:����S<g��	����j��;�U#X� ��1�<HHA84�Λ��P���5z4�W�gx{�tL?�O�X�G4��n��/Gj��X��G݈�H�9@�AA�|�͕Sw����;jx�g��g���\PTE�r�3��7��=Eiʽ[�~�����=���i��?�neY��Jͯ�O�Ι	�<1�P���5��DhW�Յ(Ѣ�˘�`��\'������21�����i�9�+b���KM���]�jNوY7�6#� �ΆR4�ۛݵA�6I���]淢�p%ф,�?�}�%2�m@˾]��^EF��&�C�'�^��(;$a�[���betu��<�ξ/M?��g��7oX�t2��y��#��O�Lc��dg�$�+D�L�K R��^P����ª i��}�8�������s/�uEq�����h����:�����I,�l�B��<ߌ�<�q&r�Qú�x�,$�\uy� အVJ�?����>E���v���]ap��X��-mS����������p
���Wa;�9~�}��f��-��i�����!�kHF��Rh��r��K�i�_`v�{�6���]�H�A�� G�a楷��:��&��<�*�^��;<��6����5�8�|�E
��?��q�l9�IxN�ē�Isy�����4!UV�M1�Ʃ�}����P66�h�����?xm��"K�Sq�;ÁV䱖H��E>#A|i~����_�n�j-�j��rX�)Ѯ���Uy�1"x����Q]טz�y�<ڤ �)g�}8�\��~��tp�:�n#�3����Jn�Ę/Ruh-ɂ�r�x0�o|S����[+��,@0���/BG>�ɔ9�1�I��<!t��-f� ����ƷF��{Rf�+�	�	�)oޗĿW��σ���X����E�6��_8��1q|g��7//����/��=7�g��H��`��d�O^�޶V~��G{]�-�2�4�_��,�錤�^h�WMm|X��զb����˱v�db0����n��m���MM��H�	F`b�X���
K`������f\3�)��u8��D��6զ�����榇�M\���k�!�eߗ�$�f��;��(�	�l���T�qb���KX&+Q�jö�ihD�ޠh���Dz�WPr�!<���<E�Ƶ����>J\#]���b����C�x�羃$Cx�8��B��|n'\�O��h�
��?����""NkhBҗ�[~�o�J�(K��*m���w�Ķ�$Y�8���)�k�}�h,�4��/��?���$���ÄQa�yq�ڶf��I�PD�t����*�uv����4RvT?�W�A�h�`?�%ǜ� P�(��T33s#��d\ۿW/��q�%Ÿ�^�y!)<>�B���t��ϧ�(n7�v�I';��a-�ur$ov��S�~�m��q�ϲ5�DrI�Yq���Č~\���b[��"�ϭH�K��B���vЅ�}76~�*�v�\�&�(�Mw�c��ǗJ.�~����:p�\�4�^, ����0U���m���Q���cF�q�R��Ӯ�D�|6ӵR��NcVP���P�5\��7P%&Д�6��5����}�w��Aww�C�e�N�iI��9��A���wS��-�畧x��hM����x|i�w�։��G_�edZ�j�x���7�h����Yf,�K���j��nn?��kO|.���it$kx��jJ��ʯF��RbѨ o(Ŗ�	m�R����\~�@a�p#��k���ro�ӽ<���1;:@H�ߋ_�Å���9����)�� 1K��l1R�ں�ē��@
�n�~Q~�M4��#�F���DL\�zЯ��J�R̓��yL�����.����!1�z\Zw��'G�|�"��Wy	1<�2D�^�����G�hpI<�]��c�T*��u�C�
ʎ̈8��s风�������c��umE��Ҧ�D)��I�L<g���#���,�2���R�����p���Ӣ�`U���r���ȕ��M�di����D�� 6���8���P��g�S����a�{���ƉZ)Wi���%��}n�j&�t���d���u\�m�#S�%a���N���٧�4����/Ѵ+HFc�zcQ.�
�I�/!�Sޠ���IQa�O}Zv����8��M~�5�)�sOL�*�֮���eN�����GNJ���ۏKö~*ћ{�K/��l�����啴7��������-��͟�-E𤎱�P�)��$�\Nh��F�6wlD@��G0ǃ���Ā'.<�X�[���Un� �?�}�	;�V���m@@���ۊD����&����2�"<+�9PK�la"a�Yk�<���;��?~V���R��?��@'x��ɕ9i�T{ᰮ̸g��^�~�O��P�-	e������0��C�7���a��q K�X���Z����
8�Ǭ�kL�w�/���	���j�x�=^�n�'1���ka|�� S�����%n���xFZ�[���D-?
���[,�e�-�ʔ!������rz��Ӕ�8Q
�i�K���:�i���:��2�ko3qF�1�i�F� ҞQi�� ��!��bC�O���k�	g�~�:^��t�M;\3:?�4�OW�A�F$( �+r0�a���?��g��.��m+M	�f4j9l��������f�g8I�7F�v�y�J�N��b%C�x���� ��I|�Ib
�ﶔg�����yL�o�;�c�L�|�:c����,(�ˡ;>�`n����b�	�O��g}�ѧ�o1�l��Z `���$�-��5�C�O)N뿚��:d�H�������ip|�k*(�qj�����z=yt3��?OM�������]H��:5��c��H�#z�H����t�����7���~,D�B�:�k4��8�1;�8�xξ��X.�"@Z�nTL?���3^s�PI��pSu��'�Q�7iT�[a�R�����z1�IM���0�B��8�'��	���+ͽ�`��yM(���{�����D��j65�:�-�
-�G�W�qR8��6��pE�:� ���R��nZ�\z�N��u*B6��f���O�z\C�: �3i�Ғ�T��5����O0�ʬ�6��2�B��l�j��	'@F Y1x�6NE�?�8��z�;��#-|���D�]#��̦�;ʝ���̮ϛ&O*�D���ŐL��3�Y�CV>��_�N�w��d�PM�L�AM�<,�s̨žr���l������)Nҏ'�8l��(C����;��g���H;�$zZ��j��za�ZWy8+������:�0�]����Z@���L��W> 8�XRK'BK�h�D����ʜ�x��%0�#��VG��t�ma�U,�k���09�a(��]�"mU�3�H�ز�pA�P����}~
ƫ�Q�/�7s�D��]��*�Ĩf�SF��w�9�p�F0�����
ȯ |v6N��n��{�����G�����ZMz��\'�֕�3E9�/eJ� "�[������ �2�c�����K���S2�Z���.�!�����4p�ei˵
�6�Ϻ}]�CeC�X�C��i-��������������G\�⭡��<3���T��7 �w:y�/}�ER��g�8�B��y�JbM�[6yK�� #v�^�#$!4���Kc�[��_s��N��8��y��e�yuN�><�<7��C��г�ljVE��A4���t��˼�R��-�}�l7�B�>�^(��G����^��ΐ�*�">��Ag-�������bT��k�A�%`���^�q����Y�<:@ b����+7��/q���ϸ���Ѱ��k��eIz;��5"_M1l�z��7�� <N	i�t5aD��-%��Jv� ?M'��K����^���S2��}:�\�6��K��;$�~���[���o{�S�@T�+�Y@�����E@x�)R��c��n*1��6��L�`iFm�Es�̮G@�����Q�D��dJ�/0�:�3B��;�L�ߨvd�1�b��j�h�����N���#���	-�e�e�ƿ$	@bx\�.O�@�܁�e{!��<��y[�d1���Q6�-j�ΡHd_< k;�<�$��I$�'"�Ɂ`QO�����t��X��I�K
���pwo&�@"XO�/�$$��$��@A�		*ٿ3a꧚2:�R��u�R��Ž0~w����[0rD��c�U�Y"�3+�E����bG���u_���2ۜ���A�f�&�q��@D �S]fvs�Gʺ����F��=c4A(f�V�j_�q���d�x$n6����q4���dI�pg�Q�!U���}2��d�D���pY�ev��cBxo)�9 wև�l��*�����a�ܶ� (�.��q�©Dz�'=�|�� �~u?<�f�u-��0��[J�D.*⟰�w�Q������+^���w{!��DL� �%���"(�U�~[1A���W9W����H��Ӝ�� ���o{bz�5�+w:
�����	!�	%�tǉ{��ǣvV�#��d�K�=M� �30�鵞j�\�{����o����Yu�r�;��1ٟ<d���lJUE�l��p<`�\I$n�Gcm�&&�Ūb�=S	�Ļ Xը��(�g]3Eݣ��+݇_[w�J�ϟ*�J���i4����E��7��:X�5��gBR��H|������B �̙�Z��#�	�X�S�~�Qȼ��+t؟X
	j��9�'��c���֤�4M�	
! ��p�ti��?W`ޟI��X^}o[pF�����D �F��l�Y��ѧ�gF̎%w���c�
�����a�	���F/�����!oη6ew$(��� ���{)�w�1�Py��;�(��5l��{�yuJ��m��h�|�R����V����O�Uk��U��&��N��JDkR�@Pg���v}�b"1~�o����b�X�l��̺�1CT��d���"�����,!� �߭�'Ё�rcVv5��t��I"&Z#�_� �_:A8��n%���N�
�硾<���8#�'V�X��uB
���+�K�|���&�#$��aaW�[v�!o��}:E�g*BvC�;�݁U����<� Q����b����"]V��?6��	��-R#�f�ȃ�xV{��������\�M�̬6^�67�4v����Z
�(��ե����� �G�B0��h���'�?,}!�%�cu o�2S9]��_`
^�q�EO'^��e]'�*�R�O6�T��l�i��?0�- �։h�&>=H�QM��m�4@�_y3���fj�95�9R�('2?�]�6!!ui	�wA�d�(�;�R����,3�"�+�	������$4z�QA�������cp�CE��CGpfKO����I�����(��!2��Nj�O76�x�CO�J���oI�8��Ć�d�bBۏȶ�C�	�����y����>
;��>�Y�a�-~������^mq6����~T�S0��mhv������m \��yo����t��'"��͹�ީ��w��>�j��b��c�,�{#܋^m��O���Tmg.��z�[�� �X�����7k��|�?NF׌	���!��1E��߭9���mGN�rݩ�'�q�gﹺv�Ã���ƃ(e����	v�����$6\��K�#TR����q�d?B^�|x;y�Ui��u�WG9B��	���A{Oh�]��L�b�F\�qV��"�q�e��p���yQ���`,�#g���Q���]��/ھ>�)Uh0�>L�ڑ��ӱG;�{�W,k ~F3)laJ�1?x��,i��hj}l瑊���c5�Rzw�F=�=��9h"��n)ۯ2�g_�C����w�����CX�,4I6"�J���qi%��E�Ǯ��z4�0u���YbE��Ot`Ty�q�o��hio"u$яȟ>��=ӵ�U�G��,*��skp�D�|�MDB���/�XHdه� �&q��M�9ԯ���O"2K �~{�Q݃7�2���Tki�}=<,s��!�~6<�xW�3v�zYG�T"�Xɗ���ẦE���WF-�8/�����Lژ��G���	�������9,3tk=A��q�|����}i�9��lþb��D��ĪZH&e/�~M�n��G:�'��Ur�`~�:���3�d:�_�- �2��.�wdT���g����@��Z�fK��Y�����V�o��Y}��ÿR�X��N�����JL{?	��V��;V�
u3}�~&�.��F�X�b҉7����k�J9��h_��| =��xgq&V��A���ftxo ��oL�E�}�"��-o;ɽ���[�oH��9�N�����~`]+ʲ�$�D�w� ��4�b%y�� ������w�*�@��{._�:m�x�?�`�dI@y����:��M'�lq��ׁu�K�?�.��@�x�6�m���U���X��m�D��g$=L�v��ѱvr&�T���d��!a[yO�<G%+p��W1�}O�-�� 0@��-khڀA�n��R�}[�
���@ �C!:���N���-���A��1���n�4H�,P�	
�>��X�HuD?�J8�Z�FoR开T@	��yq��I��3��p�%��2E���5v*I�'���k��L�+i�D�L�o�0�4k%�ƞ�ς*����Q�ͳ��$U�H0Wb5���A/�[��lB�#�'f8���'q��/|�O�8�a�WU�P�zW���֌�`��;�����GG;:�ݘ5��Աxޕo�1~z<�-F�%��\�S	�M��Ō��/�/� �+LI�B�S�N�y���w�Ӽ��z��tv;��y�ʨ�;~@n��������C�<qd�����������"-: r����Hܰ������y��U}R'_Q��^�I%�
��rG��4I=iN���M��b�X�����F� ��B��]v��
���A��OE>��OS$��j����ώ���E璂}�b��QY�,���2ѩ���^�q���8]�n�IX���0�(\vO�=���(^��a��W�ܨ�� �ZcS`����.A-���+�l^��P��߼���j�nb�^�ts( }[�gCyLG6s�q�Kؕ��Q���7�G����	������{�,�-��Ox�����U���� ��@;D���y��5�D�A�(-�t�F�*>�"hSҤc��U}�ڊ��2i��b°�>B�ڷ�_�]2�/J�e�^mX^/r��*wJ�|'%o���!��{�b]\�~��!Z;F�J�i�-r傋�ѧ�r:�l��g�7CҨ�y*?�N;e4NqB�b8׬�KTUA�*�x�ibqK�W'�ϚAYІ���~��;�����Ӆ�۰`jfbخ�?"�E��*Ɓ͙�)bb��pCg~�p�4�r�l���D'��Q@���C�a����@�B�0���P��l��]G�S�J4�B����}�T�f�P,e�o=�����'����	,��'��y^�#
@��s��=﫟��5�BR4)��>?9F�w�{���^�&��uJ^g�������ʹ������B�y����:|�'���dV�[jK�T����O*ↄ�F?+����x,Ta4��>���h�x§3�J)>p��a�6������b���s4�!2�-��'��'�Qj!�%^ �vd{�d��p��L�-�b��0|N��t�rrY�}���,�Pr��oZ��n���#\?'�����8���=G�+���l�vv��t�P���&��u����еtܱ<#���f��bOJn�g�ޤ�8_s�Vn3e)jJ��}���e$�t$���s2��ۿ[K�B���&�s���"�[�a�}�* �b�Ė�ic>��?��X�NL�L�{G�{���V²Ju����{:pk�L��Ҷ�j�hB�JN���\�E�#xok�A!�m�PZs�{�f��i&��p���΍�ꖳUj��� =,@g��Z���V�����	gh�޴xwP��a tr�� ��*;@�f��� ��.���׿z!	��!V�fy�'���e���8��#,�����sY4�h�j��~�-�T.�����l��CkV~�O׀t��}�?Ctd�L�]|,N�*3#̿����[\�~i��(d�ך;�w��+��Q�0�B�_VCuP���bj�珝�m�����/(�b8rV��o9|m������4XA!�-�f�f ΂�g�vJ��Y��]$��Q��t/��#�v��/���Mc.@r���-P���ʇٵ*���3ޱ�E
_X�B�\n$�1j[/��['QQi��z+������U8�Y)*���kA��3HV79��߲b�e�Hf���;������T�G#;�|��ç�����
%Jrڮ��P�֋) $`�B�!�R��?��V!��ܰ����)q۝�u ¡U�e@j���~�h�}3�N�0�ƻ4 :nQ]�R� ]�1D̽b��VM�QX@���y�X�CҜk�~\���0����asSw��#.T���Gq��hC�u��\�bP&`<���G@�2G~��SY�a���; `���_aơ��94��1҉������+�"ъ�.��8��=�C+����a۰�GG��Wi +I-o�Sh�Q���έ�V��"��� H�Y����齯Ĳ�cv'�h~&lc�� ��Ϧ�)j�*ydO菔ډ=֏23����K��(���v*w�TI�9f�"�yg:�G�[S=I(pF��}r�v��� ���S�u�KK����z��H^�g���
��N�=c/���&����S�G�:�ݍ�Z���L���={H��<�/��L�������z����Ć�����Z�o�3h(���"oD�3��_}�V�)3����8�>�\����r�I�.���l�8C5����5|��-��>�����Ȇ���}��� �?4C�'��ӆ�o�R=V9'b�N�h�d��;������-$/��g�BLMZ^� x�@��kνM�	0���s&s'Ilr����Z )�(Jg��gZeԗsX�n'��Z�Z��79�i�Gj�;X���>��.�E:����˲�&�i�Pz�9o����ߕP�ZV� ������-�x<��?���a�-ԇ^�&˕uV��',�o�<C �0N�i�����v4ؽg�g#�B��X�Fz���I�F���#���ځ+;8i�����Ɇ���	��OC�ef���ĸ\���b]I G$��~�y^���d������j<�(������e	��L���~�������B�!C�p�hٔC���v�1v]IɉS$��tX[�����g�t� 1_2�m���˨��Z)��W~�V���,�Ų�t����v��*D��F�́�y�F��ܒ��O/=-v�+tpH�ʤ�"\���G����gI�b�K�"5��� �;��H��o���'��aOV��&��<ކL��0Q�5����H�Rz��n±�x���mF�zW��*�j��s2�e3q
\Nʿb�#9���g��!�D��g��RmNa����`�*Y��dS<���梈�sCaB������)T�g�WGo� 4>T"�W�Nj����F�V��|�/��)s�U*��9H֊��<K�io.l��q	IOB� �$�vo 50��"wS�<aՈ+�t{:Z�^��ũ7��SBQ��;;G���ƋԨܘ9��ƞ�?��M��|�/��$ �A���/Ŕ'L�Ӑ�׷����`&�Tz�bq�KH��2}�YK
�RĽ�t��� ow*����2Mw�)�rT^ٔQ�/��VT� ��%	L9\���l�h����Pf�a�c�M=�k��e�X*_^��D2�H�z��D\�xV��[S�}��'��{4#'"2T9Rv\�m�"�S? �ʔm��;];s��Z�/��s{�ǅTt�_�޹\�Վ ܉��7s��lҘZ��QO��l0w�s��Ze���=ܟ<YP�Hªٳe���X�2⼷4�Y�n���g�a�!J�ŕJ0e )a?�7��Z�(�8H�!��F�&�mxr߹��0�F��`��ِ����z�!�d����{�muE�5.w��A,���jy���S� (M�[	�	��*K�¾�V�i�C^
��0��D�kG�&ԯ���t�ɘ<}S��w/�@)��kYd�_�,��'�hv�I��d�׆��t4('haH���F	��7����������vӒ������x��Eu���Q<�ffdi�QQ�||7-h|���-��h�˨�'��(�xh��1���s ��ma�IU)�!(�i�����whϭG��5��wȮQ���E&����>� ����P�<>`m����N>��@O�i�
���wO|���=5kTc
x�a�=�|�Q��<�E�j�>.��"%񼢞�<��@@�k�e�YeG�.C�1+f~$��"@d/���Q�Y
m�՞1U�y�^@�Yk�Q����Y�K��I3J��m�.k�A�2�0\r�:w�3 g�zS.	�Y�b�a�E-�L=�g�Rj׏���V��wA��sh&*�h�v���st�љn�:�UUP����dZ{��Q�Ȕm�)� 
"�c���a-�@D����ٞ �a~ﲙG~�n>x��Ur�P"�;`��|`��-���1���G���%E�xU=���������j���z�*p�#�q6!�nj#�E�f��1H���8�����1oC��=�܅{�;�LH(���s�,K�8�c+ BB���m�����v~|�&@���:�� ���?��.^<R:����FUE����{�$�S���6O��]�3�az#A��/2i���5�&��gt�+&F�i�=,��\%�k�a=[yG����]Ťj�=�{�4��0���Gk���w��o@{�+,@/bUގ��=����1�䠝�Ӣ�(0�����`]�
F6��.��CSO!\"���Dmz:2C��cK�`�5s���z�u@�A>���d�.���֦�>'r�ǔY�?v��9�h<�,�TE��]XU=t@����`��lj�E�ri��E�t=n����KN3��[�ʵ�ʻ���N��dF
����ޡ��Q�]�: ������CQ���J_H���Ա ���]�]�#�>��X�fFǢ�Q=�������sӑ��$<��C��9��_nO>�B��zve���)[TX��
��:$�J�X��.��9Z��ˌ�N� x�H];T���9Ab�77buw�m������F�1�	�ň�'�B�=���v�g$N���F����I���gwD�GJ=��.� j���E �M
�J��NGv��}�� ����s�GZT���)��5���پ�J���H�_�R
5���1���I�<� �ő8���BT47og�1��>��7��;������"�����g�m��O�xA�Ř���z��p?r��CX2iq��0%�gC���sF��Ԑb����l�W)�He����)��	l��@EZY���)�����>RS�\���>�#DvMt��ۦܯ��1��� "���'�@$.x�DE���'��)�jȜ�+u��<�;�j��U&�� 2TJ�>��5�]���^��z]���mO�D~-%��m��WQ�a�N��@���].�2t�	�(�#��֮>��n�Ky�P~O�gs~0F�M���8�,G�r�X~�bp��y��
�;�|�>V.1��7W��D�ABN2C��@p��?���@k��K��^GS,C8���R��Rxz"��=�;��n��	��f��)��>H��mC1݀���.�Vu�}���gG�u'���rc*�w���Fo��8��؊�#qҫ�PeZd�$9P�e�\3�Y$����O�Ϯ�1|��}	�h���MS�^)�zUg�F{i��Il�-W�h��pLF� ��V��t��c%���Y��%�U�$.H=���� ��� Yk)�N�,w���y�|,��_(fD����MY�g�0�ː�lv��^ʶ3�L�4��T��_�6�k��&�@dF5dQ�f­ɘ�H�ո&1���v�^���d����\`�"�P"=�H��uP~���f�wZkfU��cOXy�(Atrt�#7���~�#h���~"O�T�`�`u�C�Z�u�u%�m�u'��JWTo	�h���T���4Ua�ci<{S=+R^^� ��݋w1�3��0[���#�s������0K-�c�e�<�T�,#Ϙ�� ����0-��
�^ǣ ���A��������'�����DFd�`��K�fF�d� B��`�����rD���eڗ3C3ۻ]<�ɹ��'V�s�]&������U%-�	^Bfj��<�3����&��c(�&V�bs� �{<�}�Qi(P��?W��Ҭ|�W�;�b1�#���Pv��C	hzD�s� �3��sDn��֒�%=����&�-��N%~w)���#���kh^k��uJV�צ$�"l'h�*ѝS.���v8��es�1QF�~��Џӏ�nv]���2��0�R�g��ɡ�N	b"�+b�q�a�9L�N��c����{�76�c��0�( <��J(�m�������5��M0ޭ3l���tP�Lf�~㺊ݺ��5�3��e�u����I@���0��[��Y]��ᜀl��(� � (�GS��Y�K�6@3@3��>:�𘇸�g�^�8S� ~1��Q��*��iy9[�5�h#<iq�@gV�5s�81C�{*b���W�J�n�=E�
z*Yb$���R׼^��� Y�� 3S/��`M�F�}�k�+(�K�.r��^���*X�-D�Z!̣�-�8D�*��7�I�=bC��{��jZ�x����6�j�Ҝ)�}qZ �rG$�cv������T�)<�{��J"���;�X*��/=�Q�/+�1��ँ�Q�-G�^8�pv����l�c/�H�i�kK�\�{��c���H�l�/]�	�쫴tk���ׇy�";F`����2�>��QK���D,��
��~�Y�>&?���Sn��0�䛶&�$)<����ͬ��OiyBh3�Εl�h魂 T����2�S��<����% d�]k#��X4�I��:�C��X�R	��>��E����䬄S�vE� @� ��쭔�'�_Z|�*L�2n{���~�װ��Hv�UK�=y��ihz&tS:�����u�K��X=�	$Q=x�Lm~$��:t�I5+��YL+w}n�76�/ ���S,���F�b�� T(�]�����"C!z��q���O�J8ʲP�>�#4�l��4�1�H�j�ٳ��,,��Qv�Tԛ��|	I��F�:?i��䗙U���'�}�T���k*@W�ͫf�oJ�n\x�f�rC���@;& ����Z�ܗ8��}Z��ŒnHy:�hb����sΏi���+����ʼ@x�!B��OTz.1�. @��w,;�M"Z&�݈��	�b�I<r�li�.]��c�F~RtbXX��
u��)�e_�ޓ#�Eh.�"5\;#��A�B�P��4��*=}|��5g��<n�J��GΈ��f�]+僻x��&!�<ͥ�Q��w��}�m��(~Ayi���
���?IF�ꨕ���R�צ�E�z`rA�Y�ʈ.�[9R
׳c�j�}Ģ��¦E�1�8�d�d���++6��ťx�����"��^I	A�ϕ��І����u�+��C�K����V򒀅7�ʾ�J[R�7�A�KM'�΃�c�T�t�$�E�
U���<o�����+�Pj�9(��=���.�!_� e$�;��G�in}�g�Un�D���B:��&Āf;<�,��8<8�])�l�o�i���2�yF������Yd�ߐ����òK{��Tq�X�z����[Ȃ(��[�Ȝ�qeh��bŵ�|G���rG��ڟ���'ѕ9��a��3�`�����9?���:.	o��/a9\t%i�@�Q�����78��-y�_�f�?8�5)�0߭e���i�'�sf��c���ls���r;'1#W���M���J��}�{�n�.Y�zg�ƋKq<���pՔT"7T���[�j^�Ǌ�m�$���5��N3�Ȍ�ԊX��'

lg�s��^r�<>7�<-����-�0󼞯�`��� ��Mh��D��'��~���S�7fbcG����t�5�������ɹ�\׺�حx���'��r=���B���ě�D����啛��:�O���#������֪�'��;�$��*R�3�@+�4�}�12?;7J�@]Q�w��:7�L�j�f��^U8��a~���k����-�����	)��Z�T �g� =��S�d/�[���L/�e���K�i�	�&"�Du�v?�v��J��i�Vu���AlH{>,F�R5�8�#u=�薔�6²z����#F�$�[x%c�9����5B{����#�U��0(�(z���U�,��?����x��aZ���r��b��%���+3I�\��
o@���e��o� ����I%�5j�RͶx=�3�ⴊ�Rr}��4���nmj[��K.%]M�,�����mzg�?Pd��Q^85lwB}v�$ε�V}B��>'�D�uۗ��=�CHqk�!} �n�bq~�?���R([��?�d�/^���%�qn�^o�hlc�
��Do ��̽Gd��%�5���f����(J��-ml�N.8��A���%�n�I�]��5��\��|b^����R&��&��7���'��[k���T�$�.�"@����@:����(�����,L9S�w��׾��]�dhv��1�j�z����J�}p��K[[%fzX��%�O����0>/���Q3�^4�M���Qs�^�8���u�е���~�{84�N�]Ɵ(j�-!�{ڮ=�O�.Z�� D��?�k۲C�+����`�Oӳ	�����y���,n�wJ����^���9%�n��:����ME���]B7���Mh\>4|d=UػiIc2_uH��IqLv��C�{�
�w�O��OA���~��L#�At����>q3B��&�.J�k40��H:ݬ�aP���J4�r�+I�S<PBN�x�������g둏=�.�F���!W��9�Y�B�����r�ǀ�����a���c�UwI��W��3�f�Q3E��`�B�{U�<#��]v�uo�vw���!;��Kְ��-��T�W�pOPà�%�5����N0XF�|5GuhC\�c�BN�CS�L�c����+:�FvV�6�2iy +AIv�S�����$�9�q8w1
�APs(T�)^�j��\�����T���T!��/���B?i��@��s���!�X��ԥ��e^�8Z&�N�V-2?Z�K0+�.�oz�mw݊ϒ��]��%]�	�^�ή�5��ט��G��D��R��,�G9��6uD`M����"�ċ���_{h���Z�E����c��é$
E�c�=��B!T�l0��$���s!bum�+���x�ܷ+�-���a0V+�0��l"�"K��=�t��[��]���>��6��U皏i�QI-e@w�3+�?�@[�C�_�}�I���Ug�ai=-Y(��h�a�s�y�N$�j~�o��p�>����8��P];�N�}�59�	�z8��767�:��(��W���ۂC�����4&5�|�";��k+�O "�U:_k�=}�:���8�w�mB�,�Bq�q�{�<j�������$! ���
g#*Ũ5�G`����4�>3D�Xmz������э<�٭W��^m[!�ǣ+�AO3jJ�N<���N[�q6.��Y���~��I�cM`)ᄦ� �"�D���1��Q�(#C9�	��T%�	���mo�Y��Ǔ����S��q���H#j��m��t~`�X;��I�x)nc����n��@�Nو�S�&^a�����ڋjw�4I�D��OUK�[A������
~�@s�+�ֆ�J9%�ӥ-�srl���!B��h$�&Bi������th����6"aq7==
l��\�p��O( �`r��'��*V�n�	����)&4�FtT!b���U�N��L8)� �sT�5!�@0��]��~?Oq���;���b�$Fxr�<g|ħ���U׽�1�b��20D�\W����N1�eҒM���o���R��0��v��_�IW��������O|���v�3x?kE��|� �@��DzH���꣱�aF.�)����0W�2��߲!۵��\����캗��]P"U�
'�����
�
��f�����n[U�`W6*#J�8Ї��R��,RͫleE�������=�"��� �~�[�*�V�<�3�ܯ�<ϧ��c��nՋm��ݕ� �M�v�
�`2���6��@g���Pu�������(���[�x���&j��m� ��Fa��>���m�=��H<.gH�-�Ku\3ƹ?�wp O��6�jp���S:9���X}ZeW%����O!&�_n���д����B8	�
#~|V������2�g�B]y�¢(��d��\�K�%P�oh>u����%[����M�NH�J�v�V��!R�@�!�:���M�ra�#u�$�,T���¢�c%_�CU�a��hY$JR��'c7s��������)���Df�%�ڈ��75���h1 ���g4�I�x�gX��:���%���Y�-��Q��]�gTr9x��vJ����������װZ~c�N��	�����ź;���b1��i�f�r�8�0~*14�ɴ3H����$�o�� ���x�D����b�[��=��Z�f�l��� w����#�!/�(�Მ��K���d���mݽ�j��M���iM��q��`[2��s}@��s�\{j&)��dA���#��bܣX�+r�-bYL���Ct����j�����aE�a��9f�[���|�b��:sVC�Q�\-7�I� �Bm��2�d��W��R�@ Q7`�������UP��~�-�tk��7�����%����t��2�E�3_ݺ�x�D�Ĺ%���0?��2����lQ}�/�h��AFI'�";�5�p�~T�s�~7�*���(rs6.1(#�����q�}��n�Yo�F~�r*��1�K}���{��Uf�	<F�:IW��
~2��� z��#�Cf�\�k����a�v�ք۹���u��r��'���'�m̎�Վ5����a��!br��z`~.ъ�� i(p������6��$a�W�P}�w�֡�Ю bQLg�Eu	B�	z(�L�{kV����XF^���+��������Q�>��	GkՕO�-�cU%���@��C��lh�*�X�P��, HN[{� ��G2R�d�PR�/l��7Q��8A;/�~��i��a��\G�1L5�v�����(�w�̹�gy���|nN��y'�寧�����d��Ό�9������pdgc��Ȗ�R8�ڕ��Qn|�w��7U6��.��l�4�A�\�h�V��r��Q�z�S��H�iEplx��>v;l��e�\Yۓ����gL|���h����&�/�s��>�GVHEw������4�G�0�QwWJST��<�%���G� �u4s(��7c�����f�Vv�&)�-]!�Q�z/3���.,pn��Ss8$�CB������=�;�5�����Ncsh�K�YI�`���59��uJ�I�az�U\�%�=b��\�����![ĕ�vz3t�\�m y"�Q\x��|Bm��}�v�"���v�+�a4�� (߆ ~"ex�N�D>ҕ�����tDF��ULI��se�$�v& Kr����;�elU��Ńl{'�'!��C��H�|6�͙����<Q�4�T��i�
)~�YZ�c.��[��*y�����r/�ڧfi�T�#�n 4r�{�04N�����!��yI�"������(�YL��J~�A@=��<
�Uo���s=�=q����Uæ�4:��+���PK}f,L0�3O��[WȏE��ب�Bk��Y��Rn	;�}��,6ǲ��&���{\��H����h��"(�~{�t�U�ꯞ�c��06�X{�Y^uex�Y2��!y��^0�!eõ@����� ��9:�A`�8��I�MD�m�M���Ҙ�L(ifD+x��q��S�	|�m)�`sX�}DD&��˫����#2���\�!�7����/�D(�2 p_6T�J�`'�dQ��O'M�^�G4�0=yI$������X������@�L�T5�����A�N�S��������G���U����:7]hlzj���"��v�t*o����B�ɟZne�2�lc�g������ح��l������W/�i��ދ�˾%;%6�S'�ʱ���<=5�˺q�/'�-ߠ7�Fݚv�`�D���TCB0���b�G�+��Y�D��7ƌ�9�2]�5u�/�un��W[ܞ��w���P�CR�U��A_51%��`c��/�y���O�J-m00���saA�2��H�h�]T�_alu1ۍ�q���rF���:�v�8a����oIݸ���qOD�7hC���H�z!�G�8��^���fc=a+���zG��}����(���c�_iK�CSvRV$ݷ��Z�A �4q{�lw�*��& �8 �u|��Ǔݷ���"%a)��}��vø
���+�f��Z��`��d�{A��q{����\#W�m�|�H������@���|>z���H��d? �����j��6�� �ގ�hs�z��a�
�"��{�}.ݺ��s��O)xh.?�<3!���6�`��z�����bh~�F���ҺaRC�; Vh��=�٪ϞI\o��?�?��&%+8����xX��P���o	��,�q����K&��oJ�~��#~��ɾT�S.a���i��A�2����3�:8=�f�ޞ����,b6�y�9%�Pi��fF���]k�h������ۻ�]���8o%���n�����"a�p�^//7$�;����?6!�50�;PI�*�����4�p��}�b��Ŕ��0mV������m�r�� ��lsaǛ�,g���s�$�=�n\e�R�v3������'F������}������9o�/���(���}���^V$x�5M�)�1b,{;���'�+-�j�p㔰6�DZ�Js��sT���p�z~�2��>���j4��i=��X�Mr� ǌK��g������ m����`��!��?J&T��(���C�t|�g$��Z�����W� ۆZ8lL��
��p�'� @��@�=�m��ZnU�u?U[F�2~q	}�m��#A6ƅDpjղ�KO;aUP\�/`+DG�t�5R�j��CB����e���^�]J�{�����w86��T���7.��l�������F�?�)N��\gѶ���/	�x�՞*Ѫz�U�;y0�dAM(槎s���2�L�`[�:��c*$Dys��-$�h�����V�]үg:�s)0�����t8q���E\F��#y�컣(קi��	>��-`��>bfF� � *�|n��6���a�����I=.�؎L�A��ii��m��@z��]C��ȗ�#Q��Cʱ�z5��7���c{����Q��S�����*k�F˛U�ߺb[ �R�����[n`W�ٜ/�����ı6�@�^��T��1"�xU�?�߹�b
���)�4;�,m���Qv ���w�j�X$'�e<���H�\�|��΢x  �ڒlӱ_:e�(�;���[�/�ȍf�l��9�?Բ�����i �Q��"���u�S��˄�g��)��Q��|��:�s�~`��� g:�幑��aD�����`�5�?)F�# ��4�¦�j���N�`4�ݓ�T�S���W��b,��
�b�:��!��nrI���H/2�e��U��;����B��Ǉ9c�K����vS4���h����U���a$�p�r��HR=	�=_���3��K�VG3w]��WS*�U�����^>w ��aD�VX<
Ɋa{I�Ɣ#�i��,O�r��g���tQ�]G塡�?h&L�)�q �ʲZ���q����H.ad��|�~�[�ssҔ��Io'0m���&� K�;�������k�MN�*~��.euG�!fU �։:'$j{Mۗ:��Mۧ�h��I��T�di ��t>U�߈ug/}�GY~��üة�Xg��@��U&�2�C#�_z�Q�,��faɽF�/�����a��X��{B\�A�����ѪVzE��� ��D�C�n��z�6>T.�	U2%3�����:���L�& :��4������5|�ʝ�&z��OD�ܓ�ׂ��
|qTͻ��n��=Kʷ)kP��d�
dl�\NO��>4������㼊B-S_�J�Af ��u��i~[���q��}�Uu����z�0�����ױ)���w��oe�Φ/��5)"�!�|�C�;�k�"*#�I�+�NEz*�mB��15¯�f�����ӏ�šR4�ٴ��@#l&{�ݼ���L1� ՟��l��pϠ���G����V��mU�,%|*�W�� O!�8�(M3��kR]+sQc�a���/<��4�ZL&��p�YT��k�t������c����{�e
|�d޳$�胉�)v�+=!� �c�'@����Ne8ZQ�,�:A�;��� ^e��,������$5�n��Ŷ��S*�Tv��G�/a� ��vË�#�z���䌾��fA���so�~�S6�5&��&iR"��f~��z&־a��3$�Ǫ��*�b}0~l����)��3g���,����M�=�=�/ӎӡ��5���5�=]h>@����t��1`�nȡ��;��e��ҏ>u�@�B��%��c���?����
X^=f�o�J�Ȱ� �-�'K�ŷ���M"ҫ�܌� :��\���K����$c�I*���	r^�������tx��O�`%^�Y��"z���e-�Bm��"���T�D�M����yn)�S��4�4��tOºB�1��Y1��k\:7�&���V#;��O}+�)Ęv'(گR�׿�>��FE�ϒ�Ҧ��f��Y�Ax2�Beu˃��6�kF����](;����b3B��Hz���9 �`Yγ��޼\�� #��|�4(�	rJ5�y�Hl� ���NY$ݮS�l�pRn90D��ݗL����h��c���W˔'�$�$�X�S�W\ ��2���
�7�^���l��P��{��l��]%΃,�s��aЁ��� ��
{wOa!���*��Q�ݮ�L��;�8��Q$D}���}͓�����Zՠ6�4��[�0ﳧ*m�7���vJ�O,�:H��e�X��9I��jg⋴�r��P&�S^��ש��_@��C%���J;iU�t[88��'d���Y=>aJ��L��r��fˣ:�\ș�4xEn0����H��&SE�1��Q�p�H��|��Za�($��{���澝k6S�?�1o�LST2����n��2�/����i.��D�0������'=�ed��y���C�ad�c遙�	!k�$�:��n)5�_�o�(�o(����7�8��!��8Z�qeo�e�T����u��XAK)?.=*�σ����v�RE�A����l:@�L�n]�~��`�W���WY����a��-�_k��nO����/&LRp�y�G��f��K�
(�z����ǛM�l�ֶ�����C���I�b�9wy��i�[A��~��F�X����R
/G>��9� ��Q+-��	�y9sO����NYE�U���<7�F��bj������!�RA,'Df��\Tq�̧9�ٳ#����%໢��#987��N�at���sl�+�s:�	�i�$Ptk�������bB��P$m�σ,�KYR�U��(l�ji��d@���1��HHW�hW(�Ø�'��Ê�f��;�޵l��qUC����
�U� =עt����4tvU�K�8�5�Mp��3�n�L���[�7�h�R����8ŗFR>����v�֦өA��w5��o?��u���"�2�?��w$U�amF����D�XM��
J�I�F�A�v՟���&�a������9��ޢ)�pL�������/)�&��z�'r R��w�������V?�;��c"Z@����Ȫ��)��ݼ��"L�(����6��Oؓe�=~�U�S�#]"���֯h�}��*߻�/�W]_�Z��(&Ng�ɐFҜj�\7���Ӡ�Hĕ�x��j �i�R��*�ФG.����{�1Px����D��C9��fNԻ �3��c�������~����՘��(�,� ���i�N�f�;D�/��2�I�W���NbK+�Aՙ��t��c�r��z�H�h"�{�k|h��z�P��W@��J�Q?�g�$Y���q��39�I޽�:���}Mo�2��l������RH���y	�cv�JX붸ŭ;�?��/�c4�ٔ:������讨� Y���3�������	�m�JT�p����4�:�_��l0��&�U�V+Ho��zu~EÆ"@�}�.5���6��׍�p�2p!�+���Տ��hj룄�:4���dv�v;�#-_U��X�=ׯx��K#<fՏW�u瑃���:�!.�4��8��59�0����ay&����%>�*aZ)Hju��6g;#�^�+��UǶTx{D�-�u0s�!���x,[2��xq7����7�D�������i��0ӄ��͞Q��+������P��;��ӽ< � �Rl=�?��͵���i�ZЬz�6�q,������`���Cǂ	�J�b�)�t��\�R���r��;�}l�f��:�i,׉y �V��p7#d���T*cݴ���Ƙ�ҟV�&����B�	h/D�e�Ƴh&�E��|�x3��Eȍ����V(��x�}�t��j8ъ�����[�Z�$���y�� n��V�U���dޟ3ɬ4�����Q�J|0���?�3�7�����O�TZ��*	�����UT��]����S��'���8D6�xsu��V���l�@`�M`,��s�4ef&�H�&n?8ْd~�����5�l9�0�j�܎�.݇z��]�эNP$����
��Da$Z�@ϭ7ƯK�ã�F@����g�N�<K�^��I	#�#���id�m3��������+��R�Q��g�J�$Nv����4X�t���W/j��%&8N�g[r��vU�bR�u�~�ξki��HR�%��I7�8ݩGǷ��p&,��~�5�'ޫ%⏤*���K�ƺ-�r�Ds0���A���/��؀;�%+���Ԭq	�΃!U�7Z,�Y�b$s�ٔ���>�W��j�VA"<#�Z�C�Ϡ1C/`�낗ጅ��C�Au�N�C�:so �ջ���@r�)�Y���j��<�uF���T�̪�Q���*����+G�SW�k��m9r��q���+��[���}�����O�l�J{��F॓9��>����[���BL�&o5��t����~g�7�܋����SʗJ?��!��X�ю?��Af�"ĭ�Xw�,u�;w��r��we��E=�+("mLS;�ϊQ���g��AZ9$�b������0�n^�v=\�)��B�Hi�e�����ɇ<ac�q�����
�,ѾV����CIr��܈��a�9pr7���?���7q��69��(�?Mq =Xo�v����=p�*�7��f�m@{���}�-�� �^2�aɋ��D���ǬT�w?���V��vW�*b����t4�ܽ>3k�B�a�y�B���ػ:C�_c�P�߉�l�g��4��&�����(�'� ���B��D'����M�~��L��+�'��d��j%���) �@�߿��Ǉ�F�n��|���|���V!�A�5�)M��7߼���o����ȏk+��8�z�E�����t�q/I0���m���9�Lڎ�I.M@*�P����J��aix�;� aۅ�ANʙM�u$[� #�5�bT�jZ�n�<J�y�f���[�s:?�� W��@��Fl
4Ñ-��'~�\�y��u	ћ_&M%D�2M2b�"0|0��"�RE�<(s�x��%�[�ǫӖT(��{��Df�U�x3���	��?!�&��+��~rUe.�	���@�Jjw���<�e�hJ������iˈ�$t��)��o6��Q&���|�wg�f���{���)<yt�iwɼ\�7��-t1q�l����4{e��Aü����>{tk��;�R�
[�׹Q�2���5$?q��N�'�`Uc�����$b-Y�y��[���,Q���`��X���ë!yB=�٭���j����g��X���б��Cs����+Q��$���_�(�H�w�d)N�pW��-QK��<�F�W�(c؞��݌�x��J�ђ.��\��ю)��Pއ}!/W��� �����Oq�+k�R��<^���h��x:��_��,�(p�d�R���	]V+�(� >k�r��C>$e�D]��b�㘁X�s[��h7��y��`���َ�r<s�F�8)��p��Ծd31�;v�|���.0�^#��0������:�v��]�љ�?x���B �&���� W��k�5�m��K�Ŝ9ݦ��\E2����bѮ�;�"$�`�.)�,������f���#PQ{���}7���V�AUgm��Uq幋���V�)Q	�B�-���g7B����B����3֩*� �q���;�f��L'ڀ�:�n\�{�.^��3�5���ȉ:hȼ�=|/���֏z�19��Oo>�B�Wl�%6�q/��/�c='��z���:}��?����'��á6�$�GY��cY&�/��0k��[Y�no�w�O�s\)L=u�����)����,������x'���z�Zc�.FN6eU����
��n�?�|���,�s�p��S���2��J���@����[6i'UF,e���٭��8v���y�:��E���Q�P�it�j��*�ҝ֎s�'틢�����J�-���֨�R���Hŉi��sq�C�2���`EJ@�����v���]����O�k�hO0�e D�k�h���Ͽ��c�w���J�e܀�
X�6�b/q[$�����4wUC�$z���F�O0nd(��ڹy��� ��e���V�/mb����TV�F�m?��2���x¹8;>MEl����*W��[���Y���R�C���$��2�+�'�Q����A����'B)��]z��u�0�N�h^���@Fы� f��[4C���}���h �^�z�%\"��vV���D<GԂC��&�AA��p#�������4[.]�]�2�G:6+�cy9h�l�"���()bqqyE|��
4�xn&�B�;�蕣yaY��/�λp��$�߼�?�!s��.����Z��'����(�1YA�T.��v�g��23���TI	3��l����sJ�^cK�ȳ�>�U�-ja��m!��8~�J�a�7�*�ȉ,R>y��'��bX֌���~�O<4E�g;����$[h����9��Xrm	�n���]O��mm%�ǻW���rF���y���F#[���E�"mvp+�Z��Y�Yw0E��I39��+����wC�<�^��������q^%Xmn�ErF�N��a)�~j��
Q3=G��#�~:��XH��>��
P=��6�;>b�fٯ�s̋Y��1��u[�&�+�&��(DM2p`}�������
8V����g���@��ͯ��BJ~�P#�����G�
P���>_���Az�;�~��McYʅ�M��f�r�N/u��54�a�&T�.%知|BGb����(5Eq	 z�(�0�p�s��Ю9��ғP�����>���8���1�����b,P����A�\:F\��46�^��09�V*�